`timescale 1ns / 1ps


module tb_PG;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	Pattern_GeneratorA uut (
		.()
	);

	alw
	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

