`timescale 1ns/ 1ps

module Signed_Array_Multiplier_32(a, b, mul);
input [31:0] a;
input[31:0] b;
output[63:0] mul;
//Declare Wire
//Wire Partial Product
wire [31:0] pwire_0, pwire_1, pwire_2, pwire_3, pwire_4, pwire_5, pwire_6, pwire_7, pwire_8, pwire_9, pwire_10, pwire_11, pwire_12, pwire_13, pwire_14, pwire_15, pwire_16, pwire_17, pwire_18, pwire_19, pwire_20, pwire_21, pwire_22, pwire_23, pwire_24, pwire_25, pwire_26, pwire_27, pwire_28, pwire_29, pwire_30, pwire_31;
//Stage-to-Stage wire
wire [61:0] swire_1;wire [60:0] swire_2;wire [59:0] swire_3;wire [58:0] swire_4;wire [57:0] swire_5;wire [56:0] swire_6;wire [55:0] swire_7;wire [54:0] swire_8;wire [53:0] swire_9;wire [52:0] swire_10;wire [51:0] swire_11;wire [50:0] swire_12;wire [49:0] swire_13;wire [48:0] swire_14;wire [47:0] swire_15;wire [46:0] swire_16;wire [45:0] swire_17;wire [44:0] swire_18;wire [43:0] swire_19;wire [42:0] swire_20;wire [41:0] swire_21;wire [40:0] swire_22;wire [39:0] swire_23;wire [38:0] swire_24;wire [37:0] swire_25;wire [36:0] swire_26;wire [35:0] swire_27;wire [34:0] swire_28;wire [33:0] swire_29;wire [32:0] swire_30;wire [31:0] swire_31;
//Carry Propagation wire
//Stage-to-Stage wire
wire [62:0] cwire_1; wire [61:0] cwire_2; wire [60:0] cwire_3; wire [59:0] cwire_4; wire [58:0] cwire_5; wire [57:0] cwire_6; wire [56:0] cwire_7; wire [55:0] cwire_8; wire [54:0] cwire_9; wire [53:0] cwire_10; wire [52:0] cwire_11; wire [51:0] cwire_12; wire [50:0] cwire_13; wire [49:0] cwire_14; wire [48:0] cwire_15; wire [47:0] cwire_16; wire [46:0] cwire_17; wire [45:0] cwire_18; wire [44:0] cwire_19; wire [43:0] cwire_20; wire [42:0] cwire_21; wire [41:0] cwire_22; wire [40:0] cwire_23; wire [39:0] cwire_24; wire [38:0] cwire_25; wire [37:0] cwire_26; wire [36:0] cwire_27; wire [35:0] cwire_28; wire [34:0] cwire_29; wire [33:0] cwire_30; wire [32:0] cwire_31;

//Stage1 Partial Mul
ha f1(pwire_1[0], pwire_0[1], mul[1], cwire_1[0]);
fa f1_1 (pwire_1[1], pwire_0[2], cwire_1[0], swire_1[0], cwire_1[1]);
fa f1_2 (pwire_1[2], pwire_0[3], cwire_1[1], swire_1[1], cwire_1[2]);
fa f1_3 (pwire_1[3], pwire_0[4], cwire_1[2], swire_1[2], cwire_1[3]);
fa f1_4 (pwire_1[4], pwire_0[5], cwire_1[3], swire_1[3], cwire_1[4]);
fa f1_5 (pwire_1[5], pwire_0[6], cwire_1[4], swire_1[4], cwire_1[5]);
fa f1_6 (pwire_1[6], pwire_0[7], cwire_1[5], swire_1[5], cwire_1[6]);
fa f1_7 (pwire_1[7], pwire_0[8], cwire_1[6], swire_1[6], cwire_1[7]);
fa f1_8 (pwire_1[8], pwire_0[9], cwire_1[7], swire_1[7], cwire_1[8]);
fa f1_9 (pwire_1[9], pwire_0[10], cwire_1[8], swire_1[8], cwire_1[9]);
fa f1_10 (pwire_1[10], pwire_0[11], cwire_1[9], swire_1[9], cwire_1[10]);
fa f1_11 (pwire_1[11], pwire_0[12], cwire_1[10], swire_1[10], cwire_1[11]);
fa f1_12 (pwire_1[12], pwire_0[13], cwire_1[11], swire_1[11], cwire_1[12]);
fa f1_13 (pwire_1[13], pwire_0[14], cwire_1[12], swire_1[12], cwire_1[13]);
fa f1_14 (pwire_1[14], pwire_0[15], cwire_1[13], swire_1[13], cwire_1[14]);
fa f1_15 (pwire_1[15], pwire_0[16], cwire_1[14], swire_1[14], cwire_1[15]);
fa f1_16 (pwire_1[16], pwire_0[17], cwire_1[15], swire_1[15], cwire_1[16]);
fa f1_17 (pwire_1[17], pwire_0[18], cwire_1[16], swire_1[16], cwire_1[17]);
fa f1_18 (pwire_1[18], pwire_0[19], cwire_1[17], swire_1[17], cwire_1[18]);
fa f1_19 (pwire_1[19], pwire_0[20], cwire_1[18], swire_1[18], cwire_1[19]);
fa f1_20 (pwire_1[20], pwire_0[21], cwire_1[19], swire_1[19], cwire_1[20]);
fa f1_21 (pwire_1[21], pwire_0[22], cwire_1[20], swire_1[20], cwire_1[21]);
fa f1_22 (pwire_1[22], pwire_0[23], cwire_1[21], swire_1[21], cwire_1[22]);
fa f1_23 (pwire_1[23], pwire_0[24], cwire_1[22], swire_1[22], cwire_1[23]);
fa f1_24 (pwire_1[24], pwire_0[25], cwire_1[23], swire_1[23], cwire_1[24]);
fa f1_25 (pwire_1[25], pwire_0[26], cwire_1[24], swire_1[24], cwire_1[25]);
fa f1_26 (pwire_1[26], pwire_0[27], cwire_1[25], swire_1[25], cwire_1[26]);
fa f1_27 (pwire_1[27], pwire_0[28], cwire_1[26], swire_1[26], cwire_1[27]);
fa f1_28 (pwire_1[28], pwire_0[29], cwire_1[27], swire_1[27], cwire_1[28]);
fa f1_29 (pwire_1[29], pwire_0[30], cwire_1[28], swire_1[28], cwire_1[29]);
fa f1_30 (pwire_1[30], pwire_0[31], cwire_1[29], swire_1[29], cwire_1[30]);
fa f1_31 (pwire_1[31], pwire_0[31], cwire_1[30], swire_1[30], cwire_1[31]);

//Stage1Padding
fa f1__1 (pwire_1[31], pwire_0[31], cwire_1[31], swire_1[31], cwire_1[32]);
fa f1__2 (pwire_1[31], pwire_0[31], cwire_1[32], swire_1[32], cwire_1[33]);
fa f1__3 (pwire_1[31], pwire_0[31], cwire_1[33], swire_1[33], cwire_1[34]);
fa f1__4 (pwire_1[31], pwire_0[31], cwire_1[34], swire_1[34], cwire_1[35]);
fa f1__5 (pwire_1[31], pwire_0[31], cwire_1[35], swire_1[35], cwire_1[36]);
fa f1__6 (pwire_1[31], pwire_0[31], cwire_1[36], swire_1[36], cwire_1[37]);
fa f1__7 (pwire_1[31], pwire_0[31], cwire_1[37], swire_1[37], cwire_1[38]);
fa f1__8 (pwire_1[31], pwire_0[31], cwire_1[38], swire_1[38], cwire_1[39]);
fa f1__9 (pwire_1[31], pwire_0[31], cwire_1[39], swire_1[39], cwire_1[40]);
fa f1__10 (pwire_1[31], pwire_0[31], cwire_1[40], swire_1[40], cwire_1[41]);
fa f1__11 (pwire_1[31], pwire_0[31], cwire_1[41], swire_1[41], cwire_1[42]);
fa f1__12 (pwire_1[31], pwire_0[31], cwire_1[42], swire_1[42], cwire_1[43]);
fa f1__13 (pwire_1[31], pwire_0[31], cwire_1[43], swire_1[43], cwire_1[44]);
fa f1__14 (pwire_1[31], pwire_0[31], cwire_1[44], swire_1[44], cwire_1[45]);
fa f1__15 (pwire_1[31], pwire_0[31], cwire_1[45], swire_1[45], cwire_1[46]);
fa f1__16 (pwire_1[31], pwire_0[31], cwire_1[46], swire_1[46], cwire_1[47]);
fa f1__17 (pwire_1[31], pwire_0[31], cwire_1[47], swire_1[47], cwire_1[48]);
fa f1__18 (pwire_1[31], pwire_0[31], cwire_1[48], swire_1[48], cwire_1[49]);
fa f1__19 (pwire_1[31], pwire_0[31], cwire_1[49], swire_1[49], cwire_1[50]);
fa f1__20 (pwire_1[31], pwire_0[31], cwire_1[50], swire_1[50], cwire_1[51]);
fa f1__21 (pwire_1[31], pwire_0[31], cwire_1[51], swire_1[51], cwire_1[52]);
fa f1__22 (pwire_1[31], pwire_0[31], cwire_1[52], swire_1[52], cwire_1[53]);
fa f1__23 (pwire_1[31], pwire_0[31], cwire_1[53], swire_1[53], cwire_1[54]);
fa f1__24 (pwire_1[31], pwire_0[31], cwire_1[54], swire_1[54], cwire_1[55]);
fa f1__25 (pwire_1[31], pwire_0[31], cwire_1[55], swire_1[55], cwire_1[56]);
fa f1__26 (pwire_1[31], pwire_0[31], cwire_1[56], swire_1[56], cwire_1[57]);
fa f1__27 (pwire_1[31], pwire_0[31], cwire_1[57], swire_1[57], cwire_1[58]);
fa f1__28 (pwire_1[31], pwire_0[31], cwire_1[58], swire_1[58], cwire_1[59]);
fa f1__29 (pwire_1[31], pwire_0[31], cwire_1[59], swire_1[59], cwire_1[60]);
fa f1__30 (pwire_1[31], pwire_0[31], cwire_1[60], swire_1[60], cwire_1[61]);
fa f1__31 (pwire_1[31], pwire_0[31], cwire_1[61], swire_1[61], cwire_1[62]);

//Stage2 Partial Mul
ha f2(pwire_2[0], swire_1[0], mul[2], cwire_2[0]);
fa f2_1 (pwire_2[1], swire_1[1], cwire_2[0], swire_2[0], cwire_2[1]);
fa f2_2 (pwire_2[2], swire_1[2], cwire_2[1], swire_2[1], cwire_2[2]);
fa f2_3 (pwire_2[3], swire_1[3], cwire_2[2], swire_2[2], cwire_2[3]);
fa f2_4 (pwire_2[4], swire_1[4], cwire_2[3], swire_2[3], cwire_2[4]);
fa f2_5 (pwire_2[5], swire_1[5], cwire_2[4], swire_2[4], cwire_2[5]);
fa f2_6 (pwire_2[6], swire_1[6], cwire_2[5], swire_2[5], cwire_2[6]);
fa f2_7 (pwire_2[7], swire_1[7], cwire_2[6], swire_2[6], cwire_2[7]);
fa f2_8 (pwire_2[8], swire_1[8], cwire_2[7], swire_2[7], cwire_2[8]);
fa f2_9 (pwire_2[9], swire_1[9], cwire_2[8], swire_2[8], cwire_2[9]);
fa f2_10 (pwire_2[10], swire_1[10], cwire_2[9], swire_2[9], cwire_2[10]);
fa f2_11 (pwire_2[11], swire_1[11], cwire_2[10], swire_2[10], cwire_2[11]);
fa f2_12 (pwire_2[12], swire_1[12], cwire_2[11], swire_2[11], cwire_2[12]);
fa f2_13 (pwire_2[13], swire_1[13], cwire_2[12], swire_2[12], cwire_2[13]);
fa f2_14 (pwire_2[14], swire_1[14], cwire_2[13], swire_2[13], cwire_2[14]);
fa f2_15 (pwire_2[15], swire_1[15], cwire_2[14], swire_2[14], cwire_2[15]);
fa f2_16 (pwire_2[16], swire_1[16], cwire_2[15], swire_2[15], cwire_2[16]);
fa f2_17 (pwire_2[17], swire_1[17], cwire_2[16], swire_2[16], cwire_2[17]);
fa f2_18 (pwire_2[18], swire_1[18], cwire_2[17], swire_2[17], cwire_2[18]);
fa f2_19 (pwire_2[19], swire_1[19], cwire_2[18], swire_2[18], cwire_2[19]);
fa f2_20 (pwire_2[20], swire_1[20], cwire_2[19], swire_2[19], cwire_2[20]);
fa f2_21 (pwire_2[21], swire_1[21], cwire_2[20], swire_2[20], cwire_2[21]);
fa f2_22 (pwire_2[22], swire_1[22], cwire_2[21], swire_2[21], cwire_2[22]);
fa f2_23 (pwire_2[23], swire_1[23], cwire_2[22], swire_2[22], cwire_2[23]);
fa f2_24 (pwire_2[24], swire_1[24], cwire_2[23], swire_2[23], cwire_2[24]);
fa f2_25 (pwire_2[25], swire_1[25], cwire_2[24], swire_2[24], cwire_2[25]);
fa f2_26 (pwire_2[26], swire_1[26], cwire_2[25], swire_2[25], cwire_2[26]);
fa f2_27 (pwire_2[27], swire_1[27], cwire_2[26], swire_2[26], cwire_2[27]);
fa f2_28 (pwire_2[28], swire_1[28], cwire_2[27], swire_2[27], cwire_2[28]);
fa f2_29 (pwire_2[29], swire_1[29], cwire_2[28], swire_2[28], cwire_2[29]);
fa f2_30 (pwire_2[30], swire_1[30], cwire_2[29], swire_2[29], cwire_2[30]);
fa f2_31 (pwire_2[31], swire_1[31], cwire_2[30], swire_2[30], cwire_2[31]);

//Stage2Padding
fa f2__1 (pwire_2[31], swire_1[32], cwire_2[31], swire_2[31], cwire_2[32]);
fa f2__2 (pwire_2[31], swire_1[33], cwire_2[32], swire_2[32], cwire_2[33]);
fa f2__3 (pwire_2[31], swire_1[34], cwire_2[33], swire_2[33], cwire_2[34]);
fa f2__4 (pwire_2[31], swire_1[35], cwire_2[34], swire_2[34], cwire_2[35]);
fa f2__5 (pwire_2[31], swire_1[36], cwire_2[35], swire_2[35], cwire_2[36]);
fa f2__6 (pwire_2[31], swire_1[37], cwire_2[36], swire_2[36], cwire_2[37]);
fa f2__7 (pwire_2[31], swire_1[38], cwire_2[37], swire_2[37], cwire_2[38]);
fa f2__8 (pwire_2[31], swire_1[39], cwire_2[38], swire_2[38], cwire_2[39]);
fa f2__9 (pwire_2[31], swire_1[40], cwire_2[39], swire_2[39], cwire_2[40]);
fa f2__10 (pwire_2[31], swire_1[41], cwire_2[40], swire_2[40], cwire_2[41]);
fa f2__11 (pwire_2[31], swire_1[42], cwire_2[41], swire_2[41], cwire_2[42]);
fa f2__12 (pwire_2[31], swire_1[43], cwire_2[42], swire_2[42], cwire_2[43]);
fa f2__13 (pwire_2[31], swire_1[44], cwire_2[43], swire_2[43], cwire_2[44]);
fa f2__14 (pwire_2[31], swire_1[45], cwire_2[44], swire_2[44], cwire_2[45]);
fa f2__15 (pwire_2[31], swire_1[46], cwire_2[45], swire_2[45], cwire_2[46]);
fa f2__16 (pwire_2[31], swire_1[47], cwire_2[46], swire_2[46], cwire_2[47]);
fa f2__17 (pwire_2[31], swire_1[48], cwire_2[47], swire_2[47], cwire_2[48]);
fa f2__18 (pwire_2[31], swire_1[49], cwire_2[48], swire_2[48], cwire_2[49]);
fa f2__19 (pwire_2[31], swire_1[50], cwire_2[49], swire_2[49], cwire_2[50]);
fa f2__20 (pwire_2[31], swire_1[51], cwire_2[50], swire_2[50], cwire_2[51]);
fa f2__21 (pwire_2[31], swire_1[52], cwire_2[51], swire_2[51], cwire_2[52]);
fa f2__22 (pwire_2[31], swire_1[53], cwire_2[52], swire_2[52], cwire_2[53]);
fa f2__23 (pwire_2[31], swire_1[54], cwire_2[53], swire_2[53], cwire_2[54]);
fa f2__24 (pwire_2[31], swire_1[55], cwire_2[54], swire_2[54], cwire_2[55]);
fa f2__25 (pwire_2[31], swire_1[56], cwire_2[55], swire_2[55], cwire_2[56]);
fa f2__26 (pwire_2[31], swire_1[57], cwire_2[56], swire_2[56], cwire_2[57]);
fa f2__27 (pwire_2[31], swire_1[58], cwire_2[57], swire_2[57], cwire_2[58]);
fa f2__28 (pwire_2[31], swire_1[59], cwire_2[58], swire_2[58], cwire_2[59]);
fa f2__29 (pwire_2[31], swire_1[60], cwire_2[59], swire_2[59], cwire_2[60]);
fa f2__30 (pwire_2[31], swire_1[61], cwire_2[60], swire_2[60], cwire_2[61]);

//Stage3 Partial Mul
ha f3(pwire_3[0], swire_2[0], mul[3], cwire_3[0]);
fa f3_1 (pwire_3[1], swire_2[1], cwire_3[0], swire_3[0], cwire_3[1]);
fa f3_2 (pwire_3[2], swire_2[2], cwire_3[1], swire_3[1], cwire_3[2]);
fa f3_3 (pwire_3[3], swire_2[3], cwire_3[2], swire_3[2], cwire_3[3]);
fa f3_4 (pwire_3[4], swire_2[4], cwire_3[3], swire_3[3], cwire_3[4]);
fa f3_5 (pwire_3[5], swire_2[5], cwire_3[4], swire_3[4], cwire_3[5]);
fa f3_6 (pwire_3[6], swire_2[6], cwire_3[5], swire_3[5], cwire_3[6]);
fa f3_7 (pwire_3[7], swire_2[7], cwire_3[6], swire_3[6], cwire_3[7]);
fa f3_8 (pwire_3[8], swire_2[8], cwire_3[7], swire_3[7], cwire_3[8]);
fa f3_9 (pwire_3[9], swire_2[9], cwire_3[8], swire_3[8], cwire_3[9]);
fa f3_10 (pwire_3[10], swire_2[10], cwire_3[9], swire_3[9], cwire_3[10]);
fa f3_11 (pwire_3[11], swire_2[11], cwire_3[10], swire_3[10], cwire_3[11]);
fa f3_12 (pwire_3[12], swire_2[12], cwire_3[11], swire_3[11], cwire_3[12]);
fa f3_13 (pwire_3[13], swire_2[13], cwire_3[12], swire_3[12], cwire_3[13]);
fa f3_14 (pwire_3[14], swire_2[14], cwire_3[13], swire_3[13], cwire_3[14]);
fa f3_15 (pwire_3[15], swire_2[15], cwire_3[14], swire_3[14], cwire_3[15]);
fa f3_16 (pwire_3[16], swire_2[16], cwire_3[15], swire_3[15], cwire_3[16]);
fa f3_17 (pwire_3[17], swire_2[17], cwire_3[16], swire_3[16], cwire_3[17]);
fa f3_18 (pwire_3[18], swire_2[18], cwire_3[17], swire_3[17], cwire_3[18]);
fa f3_19 (pwire_3[19], swire_2[19], cwire_3[18], swire_3[18], cwire_3[19]);
fa f3_20 (pwire_3[20], swire_2[20], cwire_3[19], swire_3[19], cwire_3[20]);
fa f3_21 (pwire_3[21], swire_2[21], cwire_3[20], swire_3[20], cwire_3[21]);
fa f3_22 (pwire_3[22], swire_2[22], cwire_3[21], swire_3[21], cwire_3[22]);
fa f3_23 (pwire_3[23], swire_2[23], cwire_3[22], swire_3[22], cwire_3[23]);
fa f3_24 (pwire_3[24], swire_2[24], cwire_3[23], swire_3[23], cwire_3[24]);
fa f3_25 (pwire_3[25], swire_2[25], cwire_3[24], swire_3[24], cwire_3[25]);
fa f3_26 (pwire_3[26], swire_2[26], cwire_3[25], swire_3[25], cwire_3[26]);
fa f3_27 (pwire_3[27], swire_2[27], cwire_3[26], swire_3[26], cwire_3[27]);
fa f3_28 (pwire_3[28], swire_2[28], cwire_3[27], swire_3[27], cwire_3[28]);
fa f3_29 (pwire_3[29], swire_2[29], cwire_3[28], swire_3[28], cwire_3[29]);
fa f3_30 (pwire_3[30], swire_2[30], cwire_3[29], swire_3[29], cwire_3[30]);
fa f3_31 (pwire_3[31], swire_2[31], cwire_3[30], swire_3[30], cwire_3[31]);

//Stage3Padding
fa f3__1 (pwire_3[31], swire_2[32], cwire_3[31], swire_3[31], cwire_3[32]);
fa f3__2 (pwire_3[31], swire_2[33], cwire_3[32], swire_3[32], cwire_3[33]);
fa f3__3 (pwire_3[31], swire_2[34], cwire_3[33], swire_3[33], cwire_3[34]);
fa f3__4 (pwire_3[31], swire_2[35], cwire_3[34], swire_3[34], cwire_3[35]);
fa f3__5 (pwire_3[31], swire_2[36], cwire_3[35], swire_3[35], cwire_3[36]);
fa f3__6 (pwire_3[31], swire_2[37], cwire_3[36], swire_3[36], cwire_3[37]);
fa f3__7 (pwire_3[31], swire_2[38], cwire_3[37], swire_3[37], cwire_3[38]);
fa f3__8 (pwire_3[31], swire_2[39], cwire_3[38], swire_3[38], cwire_3[39]);
fa f3__9 (pwire_3[31], swire_2[40], cwire_3[39], swire_3[39], cwire_3[40]);
fa f3__10 (pwire_3[31], swire_2[41], cwire_3[40], swire_3[40], cwire_3[41]);
fa f3__11 (pwire_3[31], swire_2[42], cwire_3[41], swire_3[41], cwire_3[42]);
fa f3__12 (pwire_3[31], swire_2[43], cwire_3[42], swire_3[42], cwire_3[43]);
fa f3__13 (pwire_3[31], swire_2[44], cwire_3[43], swire_3[43], cwire_3[44]);
fa f3__14 (pwire_3[31], swire_2[45], cwire_3[44], swire_3[44], cwire_3[45]);
fa f3__15 (pwire_3[31], swire_2[46], cwire_3[45], swire_3[45], cwire_3[46]);
fa f3__16 (pwire_3[31], swire_2[47], cwire_3[46], swire_3[46], cwire_3[47]);
fa f3__17 (pwire_3[31], swire_2[48], cwire_3[47], swire_3[47], cwire_3[48]);
fa f3__18 (pwire_3[31], swire_2[49], cwire_3[48], swire_3[48], cwire_3[49]);
fa f3__19 (pwire_3[31], swire_2[50], cwire_3[49], swire_3[49], cwire_3[50]);
fa f3__20 (pwire_3[31], swire_2[51], cwire_3[50], swire_3[50], cwire_3[51]);
fa f3__21 (pwire_3[31], swire_2[52], cwire_3[51], swire_3[51], cwire_3[52]);
fa f3__22 (pwire_3[31], swire_2[53], cwire_3[52], swire_3[52], cwire_3[53]);
fa f3__23 (pwire_3[31], swire_2[54], cwire_3[53], swire_3[53], cwire_3[54]);
fa f3__24 (pwire_3[31], swire_2[55], cwire_3[54], swire_3[54], cwire_3[55]);
fa f3__25 (pwire_3[31], swire_2[56], cwire_3[55], swire_3[55], cwire_3[56]);
fa f3__26 (pwire_3[31], swire_2[57], cwire_3[56], swire_3[56], cwire_3[57]);
fa f3__27 (pwire_3[31], swire_2[58], cwire_3[57], swire_3[57], cwire_3[58]);
fa f3__28 (pwire_3[31], swire_2[59], cwire_3[58], swire_3[58], cwire_3[59]);
fa f3__29 (pwire_3[31], swire_2[60], cwire_3[59], swire_3[59], cwire_3[60]);

//Stage4 Partial Mul
ha f4(pwire_4[0], swire_3[0], mul[4], cwire_4[0]);
fa f4_1 (pwire_4[1], swire_3[1], cwire_4[0], swire_4[0], cwire_4[1]);
fa f4_2 (pwire_4[2], swire_3[2], cwire_4[1], swire_4[1], cwire_4[2]);
fa f4_3 (pwire_4[3], swire_3[3], cwire_4[2], swire_4[2], cwire_4[3]);
fa f4_4 (pwire_4[4], swire_3[4], cwire_4[3], swire_4[3], cwire_4[4]);
fa f4_5 (pwire_4[5], swire_3[5], cwire_4[4], swire_4[4], cwire_4[5]);
fa f4_6 (pwire_4[6], swire_3[6], cwire_4[5], swire_4[5], cwire_4[6]);
fa f4_7 (pwire_4[7], swire_3[7], cwire_4[6], swire_4[6], cwire_4[7]);
fa f4_8 (pwire_4[8], swire_3[8], cwire_4[7], swire_4[7], cwire_4[8]);
fa f4_9 (pwire_4[9], swire_3[9], cwire_4[8], swire_4[8], cwire_4[9]);
fa f4_10 (pwire_4[10], swire_3[10], cwire_4[9], swire_4[9], cwire_4[10]);
fa f4_11 (pwire_4[11], swire_3[11], cwire_4[10], swire_4[10], cwire_4[11]);
fa f4_12 (pwire_4[12], swire_3[12], cwire_4[11], swire_4[11], cwire_4[12]);
fa f4_13 (pwire_4[13], swire_3[13], cwire_4[12], swire_4[12], cwire_4[13]);
fa f4_14 (pwire_4[14], swire_3[14], cwire_4[13], swire_4[13], cwire_4[14]);
fa f4_15 (pwire_4[15], swire_3[15], cwire_4[14], swire_4[14], cwire_4[15]);
fa f4_16 (pwire_4[16], swire_3[16], cwire_4[15], swire_4[15], cwire_4[16]);
fa f4_17 (pwire_4[17], swire_3[17], cwire_4[16], swire_4[16], cwire_4[17]);
fa f4_18 (pwire_4[18], swire_3[18], cwire_4[17], swire_4[17], cwire_4[18]);
fa f4_19 (pwire_4[19], swire_3[19], cwire_4[18], swire_4[18], cwire_4[19]);
fa f4_20 (pwire_4[20], swire_3[20], cwire_4[19], swire_4[19], cwire_4[20]);
fa f4_21 (pwire_4[21], swire_3[21], cwire_4[20], swire_4[20], cwire_4[21]);
fa f4_22 (pwire_4[22], swire_3[22], cwire_4[21], swire_4[21], cwire_4[22]);
fa f4_23 (pwire_4[23], swire_3[23], cwire_4[22], swire_4[22], cwire_4[23]);
fa f4_24 (pwire_4[24], swire_3[24], cwire_4[23], swire_4[23], cwire_4[24]);
fa f4_25 (pwire_4[25], swire_3[25], cwire_4[24], swire_4[24], cwire_4[25]);
fa f4_26 (pwire_4[26], swire_3[26], cwire_4[25], swire_4[25], cwire_4[26]);
fa f4_27 (pwire_4[27], swire_3[27], cwire_4[26], swire_4[26], cwire_4[27]);
fa f4_28 (pwire_4[28], swire_3[28], cwire_4[27], swire_4[27], cwire_4[28]);
fa f4_29 (pwire_4[29], swire_3[29], cwire_4[28], swire_4[28], cwire_4[29]);
fa f4_30 (pwire_4[30], swire_3[30], cwire_4[29], swire_4[29], cwire_4[30]);
fa f4_31 (pwire_4[31], swire_3[31], cwire_4[30], swire_4[30], cwire_4[31]);

//Stage4Padding
fa f4__1 (pwire_4[31], swire_3[32], cwire_4[31], swire_4[31], cwire_4[32]);
fa f4__2 (pwire_4[31], swire_3[33], cwire_4[32], swire_4[32], cwire_4[33]);
fa f4__3 (pwire_4[31], swire_3[34], cwire_4[33], swire_4[33], cwire_4[34]);
fa f4__4 (pwire_4[31], swire_3[35], cwire_4[34], swire_4[34], cwire_4[35]);
fa f4__5 (pwire_4[31], swire_3[36], cwire_4[35], swire_4[35], cwire_4[36]);
fa f4__6 (pwire_4[31], swire_3[37], cwire_4[36], swire_4[36], cwire_4[37]);
fa f4__7 (pwire_4[31], swire_3[38], cwire_4[37], swire_4[37], cwire_4[38]);
fa f4__8 (pwire_4[31], swire_3[39], cwire_4[38], swire_4[38], cwire_4[39]);
fa f4__9 (pwire_4[31], swire_3[40], cwire_4[39], swire_4[39], cwire_4[40]);
fa f4__10 (pwire_4[31], swire_3[41], cwire_4[40], swire_4[40], cwire_4[41]);
fa f4__11 (pwire_4[31], swire_3[42], cwire_4[41], swire_4[41], cwire_4[42]);
fa f4__12 (pwire_4[31], swire_3[43], cwire_4[42], swire_4[42], cwire_4[43]);
fa f4__13 (pwire_4[31], swire_3[44], cwire_4[43], swire_4[43], cwire_4[44]);
fa f4__14 (pwire_4[31], swire_3[45], cwire_4[44], swire_4[44], cwire_4[45]);
fa f4__15 (pwire_4[31], swire_3[46], cwire_4[45], swire_4[45], cwire_4[46]);
fa f4__16 (pwire_4[31], swire_3[47], cwire_4[46], swire_4[46], cwire_4[47]);
fa f4__17 (pwire_4[31], swire_3[48], cwire_4[47], swire_4[47], cwire_4[48]);
fa f4__18 (pwire_4[31], swire_3[49], cwire_4[48], swire_4[48], cwire_4[49]);
fa f4__19 (pwire_4[31], swire_3[50], cwire_4[49], swire_4[49], cwire_4[50]);
fa f4__20 (pwire_4[31], swire_3[51], cwire_4[50], swire_4[50], cwire_4[51]);
fa f4__21 (pwire_4[31], swire_3[52], cwire_4[51], swire_4[51], cwire_4[52]);
fa f4__22 (pwire_4[31], swire_3[53], cwire_4[52], swire_4[52], cwire_4[53]);
fa f4__23 (pwire_4[31], swire_3[54], cwire_4[53], swire_4[53], cwire_4[54]);
fa f4__24 (pwire_4[31], swire_3[55], cwire_4[54], swire_4[54], cwire_4[55]);
fa f4__25 (pwire_4[31], swire_3[56], cwire_4[55], swire_4[55], cwire_4[56]);
fa f4__26 (pwire_4[31], swire_3[57], cwire_4[56], swire_4[56], cwire_4[57]);
fa f4__27 (pwire_4[31], swire_3[58], cwire_4[57], swire_4[57], cwire_4[58]);
fa f4__28 (pwire_4[31], swire_3[59], cwire_4[58], swire_4[58], cwire_4[59]);

//Stage5 Partial Mul
ha f5(pwire_5[0], swire_4[0], mul[5], cwire_5[0]);
fa f5_1 (pwire_5[1], swire_4[1], cwire_5[0], swire_5[0], cwire_5[1]);
fa f5_2 (pwire_5[2], swire_4[2], cwire_5[1], swire_5[1], cwire_5[2]);
fa f5_3 (pwire_5[3], swire_4[3], cwire_5[2], swire_5[2], cwire_5[3]);
fa f5_4 (pwire_5[4], swire_4[4], cwire_5[3], swire_5[3], cwire_5[4]);
fa f5_5 (pwire_5[5], swire_4[5], cwire_5[4], swire_5[4], cwire_5[5]);
fa f5_6 (pwire_5[6], swire_4[6], cwire_5[5], swire_5[5], cwire_5[6]);
fa f5_7 (pwire_5[7], swire_4[7], cwire_5[6], swire_5[6], cwire_5[7]);
fa f5_8 (pwire_5[8], swire_4[8], cwire_5[7], swire_5[7], cwire_5[8]);
fa f5_9 (pwire_5[9], swire_4[9], cwire_5[8], swire_5[8], cwire_5[9]);
fa f5_10 (pwire_5[10], swire_4[10], cwire_5[9], swire_5[9], cwire_5[10]);
fa f5_11 (pwire_5[11], swire_4[11], cwire_5[10], swire_5[10], cwire_5[11]);
fa f5_12 (pwire_5[12], swire_4[12], cwire_5[11], swire_5[11], cwire_5[12]);
fa f5_13 (pwire_5[13], swire_4[13], cwire_5[12], swire_5[12], cwire_5[13]);
fa f5_14 (pwire_5[14], swire_4[14], cwire_5[13], swire_5[13], cwire_5[14]);
fa f5_15 (pwire_5[15], swire_4[15], cwire_5[14], swire_5[14], cwire_5[15]);
fa f5_16 (pwire_5[16], swire_4[16], cwire_5[15], swire_5[15], cwire_5[16]);
fa f5_17 (pwire_5[17], swire_4[17], cwire_5[16], swire_5[16], cwire_5[17]);
fa f5_18 (pwire_5[18], swire_4[18], cwire_5[17], swire_5[17], cwire_5[18]);
fa f5_19 (pwire_5[19], swire_4[19], cwire_5[18], swire_5[18], cwire_5[19]);
fa f5_20 (pwire_5[20], swire_4[20], cwire_5[19], swire_5[19], cwire_5[20]);
fa f5_21 (pwire_5[21], swire_4[21], cwire_5[20], swire_5[20], cwire_5[21]);
fa f5_22 (pwire_5[22], swire_4[22], cwire_5[21], swire_5[21], cwire_5[22]);
fa f5_23 (pwire_5[23], swire_4[23], cwire_5[22], swire_5[22], cwire_5[23]);
fa f5_24 (pwire_5[24], swire_4[24], cwire_5[23], swire_5[23], cwire_5[24]);
fa f5_25 (pwire_5[25], swire_4[25], cwire_5[24], swire_5[24], cwire_5[25]);
fa f5_26 (pwire_5[26], swire_4[26], cwire_5[25], swire_5[25], cwire_5[26]);
fa f5_27 (pwire_5[27], swire_4[27], cwire_5[26], swire_5[26], cwire_5[27]);
fa f5_28 (pwire_5[28], swire_4[28], cwire_5[27], swire_5[27], cwire_5[28]);
fa f5_29 (pwire_5[29], swire_4[29], cwire_5[28], swire_5[28], cwire_5[29]);
fa f5_30 (pwire_5[30], swire_4[30], cwire_5[29], swire_5[29], cwire_5[30]);
fa f5_31 (pwire_5[31], swire_4[31], cwire_5[30], swire_5[30], cwire_5[31]);

//Stage5Padding
fa f5__1 (pwire_5[31], swire_4[32], cwire_5[31], swire_5[31], cwire_5[32]);
fa f5__2 (pwire_5[31], swire_4[33], cwire_5[32], swire_5[32], cwire_5[33]);
fa f5__3 (pwire_5[31], swire_4[34], cwire_5[33], swire_5[33], cwire_5[34]);
fa f5__4 (pwire_5[31], swire_4[35], cwire_5[34], swire_5[34], cwire_5[35]);
fa f5__5 (pwire_5[31], swire_4[36], cwire_5[35], swire_5[35], cwire_5[36]);
fa f5__6 (pwire_5[31], swire_4[37], cwire_5[36], swire_5[36], cwire_5[37]);
fa f5__7 (pwire_5[31], swire_4[38], cwire_5[37], swire_5[37], cwire_5[38]);
fa f5__8 (pwire_5[31], swire_4[39], cwire_5[38], swire_5[38], cwire_5[39]);
fa f5__9 (pwire_5[31], swire_4[40], cwire_5[39], swire_5[39], cwire_5[40]);
fa f5__10 (pwire_5[31], swire_4[41], cwire_5[40], swire_5[40], cwire_5[41]);
fa f5__11 (pwire_5[31], swire_4[42], cwire_5[41], swire_5[41], cwire_5[42]);
fa f5__12 (pwire_5[31], swire_4[43], cwire_5[42], swire_5[42], cwire_5[43]);
fa f5__13 (pwire_5[31], swire_4[44], cwire_5[43], swire_5[43], cwire_5[44]);
fa f5__14 (pwire_5[31], swire_4[45], cwire_5[44], swire_5[44], cwire_5[45]);
fa f5__15 (pwire_5[31], swire_4[46], cwire_5[45], swire_5[45], cwire_5[46]);
fa f5__16 (pwire_5[31], swire_4[47], cwire_5[46], swire_5[46], cwire_5[47]);
fa f5__17 (pwire_5[31], swire_4[48], cwire_5[47], swire_5[47], cwire_5[48]);
fa f5__18 (pwire_5[31], swire_4[49], cwire_5[48], swire_5[48], cwire_5[49]);
fa f5__19 (pwire_5[31], swire_4[50], cwire_5[49], swire_5[49], cwire_5[50]);
fa f5__20 (pwire_5[31], swire_4[51], cwire_5[50], swire_5[50], cwire_5[51]);
fa f5__21 (pwire_5[31], swire_4[52], cwire_5[51], swire_5[51], cwire_5[52]);
fa f5__22 (pwire_5[31], swire_4[53], cwire_5[52], swire_5[52], cwire_5[53]);
fa f5__23 (pwire_5[31], swire_4[54], cwire_5[53], swire_5[53], cwire_5[54]);
fa f5__24 (pwire_5[31], swire_4[55], cwire_5[54], swire_5[54], cwire_5[55]);
fa f5__25 (pwire_5[31], swire_4[56], cwire_5[55], swire_5[55], cwire_5[56]);
fa f5__26 (pwire_5[31], swire_4[57], cwire_5[56], swire_5[56], cwire_5[57]);
fa f5__27 (pwire_5[31], swire_4[58], cwire_5[57], swire_5[57], cwire_5[58]);

//Stage6 Partial Mul
ha f6(pwire_6[0], swire_5[0], mul[6], cwire_6[0]);
fa f6_1 (pwire_6[1], swire_5[1], cwire_6[0], swire_6[0], cwire_6[1]);
fa f6_2 (pwire_6[2], swire_5[2], cwire_6[1], swire_6[1], cwire_6[2]);
fa f6_3 (pwire_6[3], swire_5[3], cwire_6[2], swire_6[2], cwire_6[3]);
fa f6_4 (pwire_6[4], swire_5[4], cwire_6[3], swire_6[3], cwire_6[4]);
fa f6_5 (pwire_6[5], swire_5[5], cwire_6[4], swire_6[4], cwire_6[5]);
fa f6_6 (pwire_6[6], swire_5[6], cwire_6[5], swire_6[5], cwire_6[6]);
fa f6_7 (pwire_6[7], swire_5[7], cwire_6[6], swire_6[6], cwire_6[7]);
fa f6_8 (pwire_6[8], swire_5[8], cwire_6[7], swire_6[7], cwire_6[8]);
fa f6_9 (pwire_6[9], swire_5[9], cwire_6[8], swire_6[8], cwire_6[9]);
fa f6_10 (pwire_6[10], swire_5[10], cwire_6[9], swire_6[9], cwire_6[10]);
fa f6_11 (pwire_6[11], swire_5[11], cwire_6[10], swire_6[10], cwire_6[11]);
fa f6_12 (pwire_6[12], swire_5[12], cwire_6[11], swire_6[11], cwire_6[12]);
fa f6_13 (pwire_6[13], swire_5[13], cwire_6[12], swire_6[12], cwire_6[13]);
fa f6_14 (pwire_6[14], swire_5[14], cwire_6[13], swire_6[13], cwire_6[14]);
fa f6_15 (pwire_6[15], swire_5[15], cwire_6[14], swire_6[14], cwire_6[15]);
fa f6_16 (pwire_6[16], swire_5[16], cwire_6[15], swire_6[15], cwire_6[16]);
fa f6_17 (pwire_6[17], swire_5[17], cwire_6[16], swire_6[16], cwire_6[17]);
fa f6_18 (pwire_6[18], swire_5[18], cwire_6[17], swire_6[17], cwire_6[18]);
fa f6_19 (pwire_6[19], swire_5[19], cwire_6[18], swire_6[18], cwire_6[19]);
fa f6_20 (pwire_6[20], swire_5[20], cwire_6[19], swire_6[19], cwire_6[20]);
fa f6_21 (pwire_6[21], swire_5[21], cwire_6[20], swire_6[20], cwire_6[21]);
fa f6_22 (pwire_6[22], swire_5[22], cwire_6[21], swire_6[21], cwire_6[22]);
fa f6_23 (pwire_6[23], swire_5[23], cwire_6[22], swire_6[22], cwire_6[23]);
fa f6_24 (pwire_6[24], swire_5[24], cwire_6[23], swire_6[23], cwire_6[24]);
fa f6_25 (pwire_6[25], swire_5[25], cwire_6[24], swire_6[24], cwire_6[25]);
fa f6_26 (pwire_6[26], swire_5[26], cwire_6[25], swire_6[25], cwire_6[26]);
fa f6_27 (pwire_6[27], swire_5[27], cwire_6[26], swire_6[26], cwire_6[27]);
fa f6_28 (pwire_6[28], swire_5[28], cwire_6[27], swire_6[27], cwire_6[28]);
fa f6_29 (pwire_6[29], swire_5[29], cwire_6[28], swire_6[28], cwire_6[29]);
fa f6_30 (pwire_6[30], swire_5[30], cwire_6[29], swire_6[29], cwire_6[30]);
fa f6_31 (pwire_6[31], swire_5[31], cwire_6[30], swire_6[30], cwire_6[31]);

//Stage6Padding
fa f6__1 (pwire_6[31], swire_5[32], cwire_6[31], swire_6[31], cwire_6[32]);
fa f6__2 (pwire_6[31], swire_5[33], cwire_6[32], swire_6[32], cwire_6[33]);
fa f6__3 (pwire_6[31], swire_5[34], cwire_6[33], swire_6[33], cwire_6[34]);
fa f6__4 (pwire_6[31], swire_5[35], cwire_6[34], swire_6[34], cwire_6[35]);
fa f6__5 (pwire_6[31], swire_5[36], cwire_6[35], swire_6[35], cwire_6[36]);
fa f6__6 (pwire_6[31], swire_5[37], cwire_6[36], swire_6[36], cwire_6[37]);
fa f6__7 (pwire_6[31], swire_5[38], cwire_6[37], swire_6[37], cwire_6[38]);
fa f6__8 (pwire_6[31], swire_5[39], cwire_6[38], swire_6[38], cwire_6[39]);
fa f6__9 (pwire_6[31], swire_5[40], cwire_6[39], swire_6[39], cwire_6[40]);
fa f6__10 (pwire_6[31], swire_5[41], cwire_6[40], swire_6[40], cwire_6[41]);
fa f6__11 (pwire_6[31], swire_5[42], cwire_6[41], swire_6[41], cwire_6[42]);
fa f6__12 (pwire_6[31], swire_5[43], cwire_6[42], swire_6[42], cwire_6[43]);
fa f6__13 (pwire_6[31], swire_5[44], cwire_6[43], swire_6[43], cwire_6[44]);
fa f6__14 (pwire_6[31], swire_5[45], cwire_6[44], swire_6[44], cwire_6[45]);
fa f6__15 (pwire_6[31], swire_5[46], cwire_6[45], swire_6[45], cwire_6[46]);
fa f6__16 (pwire_6[31], swire_5[47], cwire_6[46], swire_6[46], cwire_6[47]);
fa f6__17 (pwire_6[31], swire_5[48], cwire_6[47], swire_6[47], cwire_6[48]);
fa f6__18 (pwire_6[31], swire_5[49], cwire_6[48], swire_6[48], cwire_6[49]);
fa f6__19 (pwire_6[31], swire_5[50], cwire_6[49], swire_6[49], cwire_6[50]);
fa f6__20 (pwire_6[31], swire_5[51], cwire_6[50], swire_6[50], cwire_6[51]);
fa f6__21 (pwire_6[31], swire_5[52], cwire_6[51], swire_6[51], cwire_6[52]);
fa f6__22 (pwire_6[31], swire_5[53], cwire_6[52], swire_6[52], cwire_6[53]);
fa f6__23 (pwire_6[31], swire_5[54], cwire_6[53], swire_6[53], cwire_6[54]);
fa f6__24 (pwire_6[31], swire_5[55], cwire_6[54], swire_6[54], cwire_6[55]);
fa f6__25 (pwire_6[31], swire_5[56], cwire_6[55], swire_6[55], cwire_6[56]);
fa f6__26 (pwire_6[31], swire_5[57], cwire_6[56], swire_6[56], cwire_6[57]);

//Stage7 Partial Mul
ha f7(pwire_7[0], swire_6[0], mul[7], cwire_7[0]);
fa f7_1 (pwire_7[1], swire_6[1], cwire_7[0], swire_7[0], cwire_7[1]);
fa f7_2 (pwire_7[2], swire_6[2], cwire_7[1], swire_7[1], cwire_7[2]);
fa f7_3 (pwire_7[3], swire_6[3], cwire_7[2], swire_7[2], cwire_7[3]);
fa f7_4 (pwire_7[4], swire_6[4], cwire_7[3], swire_7[3], cwire_7[4]);
fa f7_5 (pwire_7[5], swire_6[5], cwire_7[4], swire_7[4], cwire_7[5]);
fa f7_6 (pwire_7[6], swire_6[6], cwire_7[5], swire_7[5], cwire_7[6]);
fa f7_7 (pwire_7[7], swire_6[7], cwire_7[6], swire_7[6], cwire_7[7]);
fa f7_8 (pwire_7[8], swire_6[8], cwire_7[7], swire_7[7], cwire_7[8]);
fa f7_9 (pwire_7[9], swire_6[9], cwire_7[8], swire_7[8], cwire_7[9]);
fa f7_10 (pwire_7[10], swire_6[10], cwire_7[9], swire_7[9], cwire_7[10]);
fa f7_11 (pwire_7[11], swire_6[11], cwire_7[10], swire_7[10], cwire_7[11]);
fa f7_12 (pwire_7[12], swire_6[12], cwire_7[11], swire_7[11], cwire_7[12]);
fa f7_13 (pwire_7[13], swire_6[13], cwire_7[12], swire_7[12], cwire_7[13]);
fa f7_14 (pwire_7[14], swire_6[14], cwire_7[13], swire_7[13], cwire_7[14]);
fa f7_15 (pwire_7[15], swire_6[15], cwire_7[14], swire_7[14], cwire_7[15]);
fa f7_16 (pwire_7[16], swire_6[16], cwire_7[15], swire_7[15], cwire_7[16]);
fa f7_17 (pwire_7[17], swire_6[17], cwire_7[16], swire_7[16], cwire_7[17]);
fa f7_18 (pwire_7[18], swire_6[18], cwire_7[17], swire_7[17], cwire_7[18]);
fa f7_19 (pwire_7[19], swire_6[19], cwire_7[18], swire_7[18], cwire_7[19]);
fa f7_20 (pwire_7[20], swire_6[20], cwire_7[19], swire_7[19], cwire_7[20]);
fa f7_21 (pwire_7[21], swire_6[21], cwire_7[20], swire_7[20], cwire_7[21]);
fa f7_22 (pwire_7[22], swire_6[22], cwire_7[21], swire_7[21], cwire_7[22]);
fa f7_23 (pwire_7[23], swire_6[23], cwire_7[22], swire_7[22], cwire_7[23]);
fa f7_24 (pwire_7[24], swire_6[24], cwire_7[23], swire_7[23], cwire_7[24]);
fa f7_25 (pwire_7[25], swire_6[25], cwire_7[24], swire_7[24], cwire_7[25]);
fa f7_26 (pwire_7[26], swire_6[26], cwire_7[25], swire_7[25], cwire_7[26]);
fa f7_27 (pwire_7[27], swire_6[27], cwire_7[26], swire_7[26], cwire_7[27]);
fa f7_28 (pwire_7[28], swire_6[28], cwire_7[27], swire_7[27], cwire_7[28]);
fa f7_29 (pwire_7[29], swire_6[29], cwire_7[28], swire_7[28], cwire_7[29]);
fa f7_30 (pwire_7[30], swire_6[30], cwire_7[29], swire_7[29], cwire_7[30]);
fa f7_31 (pwire_7[31], swire_6[31], cwire_7[30], swire_7[30], cwire_7[31]);

//Stage7Padding
fa f7__1 (pwire_7[31], swire_6[32], cwire_7[31], swire_7[31], cwire_7[32]);
fa f7__2 (pwire_7[31], swire_6[33], cwire_7[32], swire_7[32], cwire_7[33]);
fa f7__3 (pwire_7[31], swire_6[34], cwire_7[33], swire_7[33], cwire_7[34]);
fa f7__4 (pwire_7[31], swire_6[35], cwire_7[34], swire_7[34], cwire_7[35]);
fa f7__5 (pwire_7[31], swire_6[36], cwire_7[35], swire_7[35], cwire_7[36]);
fa f7__6 (pwire_7[31], swire_6[37], cwire_7[36], swire_7[36], cwire_7[37]);
fa f7__7 (pwire_7[31], swire_6[38], cwire_7[37], swire_7[37], cwire_7[38]);
fa f7__8 (pwire_7[31], swire_6[39], cwire_7[38], swire_7[38], cwire_7[39]);
fa f7__9 (pwire_7[31], swire_6[40], cwire_7[39], swire_7[39], cwire_7[40]);
fa f7__10 (pwire_7[31], swire_6[41], cwire_7[40], swire_7[40], cwire_7[41]);
fa f7__11 (pwire_7[31], swire_6[42], cwire_7[41], swire_7[41], cwire_7[42]);
fa f7__12 (pwire_7[31], swire_6[43], cwire_7[42], swire_7[42], cwire_7[43]);
fa f7__13 (pwire_7[31], swire_6[44], cwire_7[43], swire_7[43], cwire_7[44]);
fa f7__14 (pwire_7[31], swire_6[45], cwire_7[44], swire_7[44], cwire_7[45]);
fa f7__15 (pwire_7[31], swire_6[46], cwire_7[45], swire_7[45], cwire_7[46]);
fa f7__16 (pwire_7[31], swire_6[47], cwire_7[46], swire_7[46], cwire_7[47]);
fa f7__17 (pwire_7[31], swire_6[48], cwire_7[47], swire_7[47], cwire_7[48]);
fa f7__18 (pwire_7[31], swire_6[49], cwire_7[48], swire_7[48], cwire_7[49]);
fa f7__19 (pwire_7[31], swire_6[50], cwire_7[49], swire_7[49], cwire_7[50]);
fa f7__20 (pwire_7[31], swire_6[51], cwire_7[50], swire_7[50], cwire_7[51]);
fa f7__21 (pwire_7[31], swire_6[52], cwire_7[51], swire_7[51], cwire_7[52]);
fa f7__22 (pwire_7[31], swire_6[53], cwire_7[52], swire_7[52], cwire_7[53]);
fa f7__23 (pwire_7[31], swire_6[54], cwire_7[53], swire_7[53], cwire_7[54]);
fa f7__24 (pwire_7[31], swire_6[55], cwire_7[54], swire_7[54], cwire_7[55]);
fa f7__25 (pwire_7[31], swire_6[56], cwire_7[55], swire_7[55], cwire_7[56]);

//Stage8 Partial Mul
ha f8(pwire_8[0], swire_7[0], mul[8], cwire_8[0]);
fa f8_1 (pwire_8[1], swire_7[1], cwire_8[0], swire_8[0], cwire_8[1]);
fa f8_2 (pwire_8[2], swire_7[2], cwire_8[1], swire_8[1], cwire_8[2]);
fa f8_3 (pwire_8[3], swire_7[3], cwire_8[2], swire_8[2], cwire_8[3]);
fa f8_4 (pwire_8[4], swire_7[4], cwire_8[3], swire_8[3], cwire_8[4]);
fa f8_5 (pwire_8[5], swire_7[5], cwire_8[4], swire_8[4], cwire_8[5]);
fa f8_6 (pwire_8[6], swire_7[6], cwire_8[5], swire_8[5], cwire_8[6]);
fa f8_7 (pwire_8[7], swire_7[7], cwire_8[6], swire_8[6], cwire_8[7]);
fa f8_8 (pwire_8[8], swire_7[8], cwire_8[7], swire_8[7], cwire_8[8]);
fa f8_9 (pwire_8[9], swire_7[9], cwire_8[8], swire_8[8], cwire_8[9]);
fa f8_10 (pwire_8[10], swire_7[10], cwire_8[9], swire_8[9], cwire_8[10]);
fa f8_11 (pwire_8[11], swire_7[11], cwire_8[10], swire_8[10], cwire_8[11]);
fa f8_12 (pwire_8[12], swire_7[12], cwire_8[11], swire_8[11], cwire_8[12]);
fa f8_13 (pwire_8[13], swire_7[13], cwire_8[12], swire_8[12], cwire_8[13]);
fa f8_14 (pwire_8[14], swire_7[14], cwire_8[13], swire_8[13], cwire_8[14]);
fa f8_15 (pwire_8[15], swire_7[15], cwire_8[14], swire_8[14], cwire_8[15]);
fa f8_16 (pwire_8[16], swire_7[16], cwire_8[15], swire_8[15], cwire_8[16]);
fa f8_17 (pwire_8[17], swire_7[17], cwire_8[16], swire_8[16], cwire_8[17]);
fa f8_18 (pwire_8[18], swire_7[18], cwire_8[17], swire_8[17], cwire_8[18]);
fa f8_19 (pwire_8[19], swire_7[19], cwire_8[18], swire_8[18], cwire_8[19]);
fa f8_20 (pwire_8[20], swire_7[20], cwire_8[19], swire_8[19], cwire_8[20]);
fa f8_21 (pwire_8[21], swire_7[21], cwire_8[20], swire_8[20], cwire_8[21]);
fa f8_22 (pwire_8[22], swire_7[22], cwire_8[21], swire_8[21], cwire_8[22]);
fa f8_23 (pwire_8[23], swire_7[23], cwire_8[22], swire_8[22], cwire_8[23]);
fa f8_24 (pwire_8[24], swire_7[24], cwire_8[23], swire_8[23], cwire_8[24]);
fa f8_25 (pwire_8[25], swire_7[25], cwire_8[24], swire_8[24], cwire_8[25]);
fa f8_26 (pwire_8[26], swire_7[26], cwire_8[25], swire_8[25], cwire_8[26]);
fa f8_27 (pwire_8[27], swire_7[27], cwire_8[26], swire_8[26], cwire_8[27]);
fa f8_28 (pwire_8[28], swire_7[28], cwire_8[27], swire_8[27], cwire_8[28]);
fa f8_29 (pwire_8[29], swire_7[29], cwire_8[28], swire_8[28], cwire_8[29]);
fa f8_30 (pwire_8[30], swire_7[30], cwire_8[29], swire_8[29], cwire_8[30]);
fa f8_31 (pwire_8[31], swire_7[31], cwire_8[30], swire_8[30], cwire_8[31]);

//Stage8Padding
fa f8__1 (pwire_8[31], swire_7[32], cwire_8[31], swire_8[31], cwire_8[32]);
fa f8__2 (pwire_8[31], swire_7[33], cwire_8[32], swire_8[32], cwire_8[33]);
fa f8__3 (pwire_8[31], swire_7[34], cwire_8[33], swire_8[33], cwire_8[34]);
fa f8__4 (pwire_8[31], swire_7[35], cwire_8[34], swire_8[34], cwire_8[35]);
fa f8__5 (pwire_8[31], swire_7[36], cwire_8[35], swire_8[35], cwire_8[36]);
fa f8__6 (pwire_8[31], swire_7[37], cwire_8[36], swire_8[36], cwire_8[37]);
fa f8__7 (pwire_8[31], swire_7[38], cwire_8[37], swire_8[37], cwire_8[38]);
fa f8__8 (pwire_8[31], swire_7[39], cwire_8[38], swire_8[38], cwire_8[39]);
fa f8__9 (pwire_8[31], swire_7[40], cwire_8[39], swire_8[39], cwire_8[40]);
fa f8__10 (pwire_8[31], swire_7[41], cwire_8[40], swire_8[40], cwire_8[41]);
fa f8__11 (pwire_8[31], swire_7[42], cwire_8[41], swire_8[41], cwire_8[42]);
fa f8__12 (pwire_8[31], swire_7[43], cwire_8[42], swire_8[42], cwire_8[43]);
fa f8__13 (pwire_8[31], swire_7[44], cwire_8[43], swire_8[43], cwire_8[44]);
fa f8__14 (pwire_8[31], swire_7[45], cwire_8[44], swire_8[44], cwire_8[45]);
fa f8__15 (pwire_8[31], swire_7[46], cwire_8[45], swire_8[45], cwire_8[46]);
fa f8__16 (pwire_8[31], swire_7[47], cwire_8[46], swire_8[46], cwire_8[47]);
fa f8__17 (pwire_8[31], swire_7[48], cwire_8[47], swire_8[47], cwire_8[48]);
fa f8__18 (pwire_8[31], swire_7[49], cwire_8[48], swire_8[48], cwire_8[49]);
fa f8__19 (pwire_8[31], swire_7[50], cwire_8[49], swire_8[49], cwire_8[50]);
fa f8__20 (pwire_8[31], swire_7[51], cwire_8[50], swire_8[50], cwire_8[51]);
fa f8__21 (pwire_8[31], swire_7[52], cwire_8[51], swire_8[51], cwire_8[52]);
fa f8__22 (pwire_8[31], swire_7[53], cwire_8[52], swire_8[52], cwire_8[53]);
fa f8__23 (pwire_8[31], swire_7[54], cwire_8[53], swire_8[53], cwire_8[54]);
fa f8__24 (pwire_8[31], swire_7[55], cwire_8[54], swire_8[54], cwire_8[55]);

//Stage9 Partial Mul
ha f9(pwire_9[0], swire_8[0], mul[9], cwire_9[0]);
fa f9_1 (pwire_9[1], swire_8[1], cwire_9[0], swire_9[0], cwire_9[1]);
fa f9_2 (pwire_9[2], swire_8[2], cwire_9[1], swire_9[1], cwire_9[2]);
fa f9_3 (pwire_9[3], swire_8[3], cwire_9[2], swire_9[2], cwire_9[3]);
fa f9_4 (pwire_9[4], swire_8[4], cwire_9[3], swire_9[3], cwire_9[4]);
fa f9_5 (pwire_9[5], swire_8[5], cwire_9[4], swire_9[4], cwire_9[5]);
fa f9_6 (pwire_9[6], swire_8[6], cwire_9[5], swire_9[5], cwire_9[6]);
fa f9_7 (pwire_9[7], swire_8[7], cwire_9[6], swire_9[6], cwire_9[7]);
fa f9_8 (pwire_9[8], swire_8[8], cwire_9[7], swire_9[7], cwire_9[8]);
fa f9_9 (pwire_9[9], swire_8[9], cwire_9[8], swire_9[8], cwire_9[9]);
fa f9_10 (pwire_9[10], swire_8[10], cwire_9[9], swire_9[9], cwire_9[10]);
fa f9_11 (pwire_9[11], swire_8[11], cwire_9[10], swire_9[10], cwire_9[11]);
fa f9_12 (pwire_9[12], swire_8[12], cwire_9[11], swire_9[11], cwire_9[12]);
fa f9_13 (pwire_9[13], swire_8[13], cwire_9[12], swire_9[12], cwire_9[13]);
fa f9_14 (pwire_9[14], swire_8[14], cwire_9[13], swire_9[13], cwire_9[14]);
fa f9_15 (pwire_9[15], swire_8[15], cwire_9[14], swire_9[14], cwire_9[15]);
fa f9_16 (pwire_9[16], swire_8[16], cwire_9[15], swire_9[15], cwire_9[16]);
fa f9_17 (pwire_9[17], swire_8[17], cwire_9[16], swire_9[16], cwire_9[17]);
fa f9_18 (pwire_9[18], swire_8[18], cwire_9[17], swire_9[17], cwire_9[18]);
fa f9_19 (pwire_9[19], swire_8[19], cwire_9[18], swire_9[18], cwire_9[19]);
fa f9_20 (pwire_9[20], swire_8[20], cwire_9[19], swire_9[19], cwire_9[20]);
fa f9_21 (pwire_9[21], swire_8[21], cwire_9[20], swire_9[20], cwire_9[21]);
fa f9_22 (pwire_9[22], swire_8[22], cwire_9[21], swire_9[21], cwire_9[22]);
fa f9_23 (pwire_9[23], swire_8[23], cwire_9[22], swire_9[22], cwire_9[23]);
fa f9_24 (pwire_9[24], swire_8[24], cwire_9[23], swire_9[23], cwire_9[24]);
fa f9_25 (pwire_9[25], swire_8[25], cwire_9[24], swire_9[24], cwire_9[25]);
fa f9_26 (pwire_9[26], swire_8[26], cwire_9[25], swire_9[25], cwire_9[26]);
fa f9_27 (pwire_9[27], swire_8[27], cwire_9[26], swire_9[26], cwire_9[27]);
fa f9_28 (pwire_9[28], swire_8[28], cwire_9[27], swire_9[27], cwire_9[28]);
fa f9_29 (pwire_9[29], swire_8[29], cwire_9[28], swire_9[28], cwire_9[29]);
fa f9_30 (pwire_9[30], swire_8[30], cwire_9[29], swire_9[29], cwire_9[30]);
fa f9_31 (pwire_9[31], swire_8[31], cwire_9[30], swire_9[30], cwire_9[31]);

//Stage9Padding
fa f9__1 (pwire_9[31], swire_8[32], cwire_9[31], swire_9[31], cwire_9[32]);
fa f9__2 (pwire_9[31], swire_8[33], cwire_9[32], swire_9[32], cwire_9[33]);
fa f9__3 (pwire_9[31], swire_8[34], cwire_9[33], swire_9[33], cwire_9[34]);
fa f9__4 (pwire_9[31], swire_8[35], cwire_9[34], swire_9[34], cwire_9[35]);
fa f9__5 (pwire_9[31], swire_8[36], cwire_9[35], swire_9[35], cwire_9[36]);
fa f9__6 (pwire_9[31], swire_8[37], cwire_9[36], swire_9[36], cwire_9[37]);
fa f9__7 (pwire_9[31], swire_8[38], cwire_9[37], swire_9[37], cwire_9[38]);
fa f9__8 (pwire_9[31], swire_8[39], cwire_9[38], swire_9[38], cwire_9[39]);
fa f9__9 (pwire_9[31], swire_8[40], cwire_9[39], swire_9[39], cwire_9[40]);
fa f9__10 (pwire_9[31], swire_8[41], cwire_9[40], swire_9[40], cwire_9[41]);
fa f9__11 (pwire_9[31], swire_8[42], cwire_9[41], swire_9[41], cwire_9[42]);
fa f9__12 (pwire_9[31], swire_8[43], cwire_9[42], swire_9[42], cwire_9[43]);
fa f9__13 (pwire_9[31], swire_8[44], cwire_9[43], swire_9[43], cwire_9[44]);
fa f9__14 (pwire_9[31], swire_8[45], cwire_9[44], swire_9[44], cwire_9[45]);
fa f9__15 (pwire_9[31], swire_8[46], cwire_9[45], swire_9[45], cwire_9[46]);
fa f9__16 (pwire_9[31], swire_8[47], cwire_9[46], swire_9[46], cwire_9[47]);
fa f9__17 (pwire_9[31], swire_8[48], cwire_9[47], swire_9[47], cwire_9[48]);
fa f9__18 (pwire_9[31], swire_8[49], cwire_9[48], swire_9[48], cwire_9[49]);
fa f9__19 (pwire_9[31], swire_8[50], cwire_9[49], swire_9[49], cwire_9[50]);
fa f9__20 (pwire_9[31], swire_8[51], cwire_9[50], swire_9[50], cwire_9[51]);
fa f9__21 (pwire_9[31], swire_8[52], cwire_9[51], swire_9[51], cwire_9[52]);
fa f9__22 (pwire_9[31], swire_8[53], cwire_9[52], swire_9[52], cwire_9[53]);
fa f9__23 (pwire_9[31], swire_8[54], cwire_9[53], swire_9[53], cwire_9[54]);

//Stage10 Partial Mul
ha f10(pwire_10[0], swire_9[0], mul[10], cwire_10[0]);
fa f10_1 (pwire_10[1], swire_9[1], cwire_10[0], swire_10[0], cwire_10[1]);
fa f10_2 (pwire_10[2], swire_9[2], cwire_10[1], swire_10[1], cwire_10[2]);
fa f10_3 (pwire_10[3], swire_9[3], cwire_10[2], swire_10[2], cwire_10[3]);
fa f10_4 (pwire_10[4], swire_9[4], cwire_10[3], swire_10[3], cwire_10[4]);
fa f10_5 (pwire_10[5], swire_9[5], cwire_10[4], swire_10[4], cwire_10[5]);
fa f10_6 (pwire_10[6], swire_9[6], cwire_10[5], swire_10[5], cwire_10[6]);
fa f10_7 (pwire_10[7], swire_9[7], cwire_10[6], swire_10[6], cwire_10[7]);
fa f10_8 (pwire_10[8], swire_9[8], cwire_10[7], swire_10[7], cwire_10[8]);
fa f10_9 (pwire_10[9], swire_9[9], cwire_10[8], swire_10[8], cwire_10[9]);
fa f10_10 (pwire_10[10], swire_9[10], cwire_10[9], swire_10[9], cwire_10[10]);
fa f10_11 (pwire_10[11], swire_9[11], cwire_10[10], swire_10[10], cwire_10[11]);
fa f10_12 (pwire_10[12], swire_9[12], cwire_10[11], swire_10[11], cwire_10[12]);
fa f10_13 (pwire_10[13], swire_9[13], cwire_10[12], swire_10[12], cwire_10[13]);
fa f10_14 (pwire_10[14], swire_9[14], cwire_10[13], swire_10[13], cwire_10[14]);
fa f10_15 (pwire_10[15], swire_9[15], cwire_10[14], swire_10[14], cwire_10[15]);
fa f10_16 (pwire_10[16], swire_9[16], cwire_10[15], swire_10[15], cwire_10[16]);
fa f10_17 (pwire_10[17], swire_9[17], cwire_10[16], swire_10[16], cwire_10[17]);
fa f10_18 (pwire_10[18], swire_9[18], cwire_10[17], swire_10[17], cwire_10[18]);
fa f10_19 (pwire_10[19], swire_9[19], cwire_10[18], swire_10[18], cwire_10[19]);
fa f10_20 (pwire_10[20], swire_9[20], cwire_10[19], swire_10[19], cwire_10[20]);
fa f10_21 (pwire_10[21], swire_9[21], cwire_10[20], swire_10[20], cwire_10[21]);
fa f10_22 (pwire_10[22], swire_9[22], cwire_10[21], swire_10[21], cwire_10[22]);
fa f10_23 (pwire_10[23], swire_9[23], cwire_10[22], swire_10[22], cwire_10[23]);
fa f10_24 (pwire_10[24], swire_9[24], cwire_10[23], swire_10[23], cwire_10[24]);
fa f10_25 (pwire_10[25], swire_9[25], cwire_10[24], swire_10[24], cwire_10[25]);
fa f10_26 (pwire_10[26], swire_9[26], cwire_10[25], swire_10[25], cwire_10[26]);
fa f10_27 (pwire_10[27], swire_9[27], cwire_10[26], swire_10[26], cwire_10[27]);
fa f10_28 (pwire_10[28], swire_9[28], cwire_10[27], swire_10[27], cwire_10[28]);
fa f10_29 (pwire_10[29], swire_9[29], cwire_10[28], swire_10[28], cwire_10[29]);
fa f10_30 (pwire_10[30], swire_9[30], cwire_10[29], swire_10[29], cwire_10[30]);
fa f10_31 (pwire_10[31], swire_9[31], cwire_10[30], swire_10[30], cwire_10[31]);

//Stage10Padding
fa f10__1 (pwire_10[31], swire_9[32], cwire_10[31], swire_10[31], cwire_10[32]);
fa f10__2 (pwire_10[31], swire_9[33], cwire_10[32], swire_10[32], cwire_10[33]);
fa f10__3 (pwire_10[31], swire_9[34], cwire_10[33], swire_10[33], cwire_10[34]);
fa f10__4 (pwire_10[31], swire_9[35], cwire_10[34], swire_10[34], cwire_10[35]);
fa f10__5 (pwire_10[31], swire_9[36], cwire_10[35], swire_10[35], cwire_10[36]);
fa f10__6 (pwire_10[31], swire_9[37], cwire_10[36], swire_10[36], cwire_10[37]);
fa f10__7 (pwire_10[31], swire_9[38], cwire_10[37], swire_10[37], cwire_10[38]);
fa f10__8 (pwire_10[31], swire_9[39], cwire_10[38], swire_10[38], cwire_10[39]);
fa f10__9 (pwire_10[31], swire_9[40], cwire_10[39], swire_10[39], cwire_10[40]);
fa f10__10 (pwire_10[31], swire_9[41], cwire_10[40], swire_10[40], cwire_10[41]);
fa f10__11 (pwire_10[31], swire_9[42], cwire_10[41], swire_10[41], cwire_10[42]);
fa f10__12 (pwire_10[31], swire_9[43], cwire_10[42], swire_10[42], cwire_10[43]);
fa f10__13 (pwire_10[31], swire_9[44], cwire_10[43], swire_10[43], cwire_10[44]);
fa f10__14 (pwire_10[31], swire_9[45], cwire_10[44], swire_10[44], cwire_10[45]);
fa f10__15 (pwire_10[31], swire_9[46], cwire_10[45], swire_10[45], cwire_10[46]);
fa f10__16 (pwire_10[31], swire_9[47], cwire_10[46], swire_10[46], cwire_10[47]);
fa f10__17 (pwire_10[31], swire_9[48], cwire_10[47], swire_10[47], cwire_10[48]);
fa f10__18 (pwire_10[31], swire_9[49], cwire_10[48], swire_10[48], cwire_10[49]);
fa f10__19 (pwire_10[31], swire_9[50], cwire_10[49], swire_10[49], cwire_10[50]);
fa f10__20 (pwire_10[31], swire_9[51], cwire_10[50], swire_10[50], cwire_10[51]);
fa f10__21 (pwire_10[31], swire_9[52], cwire_10[51], swire_10[51], cwire_10[52]);
fa f10__22 (pwire_10[31], swire_9[53], cwire_10[52], swire_10[52], cwire_10[53]);

//Stage11 Partial Mul
ha f11(pwire_11[0], swire_10[0], mul[11], cwire_11[0]);
fa f11_1 (pwire_11[1], swire_10[1], cwire_11[0], swire_11[0], cwire_11[1]);
fa f11_2 (pwire_11[2], swire_10[2], cwire_11[1], swire_11[1], cwire_11[2]);
fa f11_3 (pwire_11[3], swire_10[3], cwire_11[2], swire_11[2], cwire_11[3]);
fa f11_4 (pwire_11[4], swire_10[4], cwire_11[3], swire_11[3], cwire_11[4]);
fa f11_5 (pwire_11[5], swire_10[5], cwire_11[4], swire_11[4], cwire_11[5]);
fa f11_6 (pwire_11[6], swire_10[6], cwire_11[5], swire_11[5], cwire_11[6]);
fa f11_7 (pwire_11[7], swire_10[7], cwire_11[6], swire_11[6], cwire_11[7]);
fa f11_8 (pwire_11[8], swire_10[8], cwire_11[7], swire_11[7], cwire_11[8]);
fa f11_9 (pwire_11[9], swire_10[9], cwire_11[8], swire_11[8], cwire_11[9]);
fa f11_10 (pwire_11[10], swire_10[10], cwire_11[9], swire_11[9], cwire_11[10]);
fa f11_11 (pwire_11[11], swire_10[11], cwire_11[10], swire_11[10], cwire_11[11]);
fa f11_12 (pwire_11[12], swire_10[12], cwire_11[11], swire_11[11], cwire_11[12]);
fa f11_13 (pwire_11[13], swire_10[13], cwire_11[12], swire_11[12], cwire_11[13]);
fa f11_14 (pwire_11[14], swire_10[14], cwire_11[13], swire_11[13], cwire_11[14]);
fa f11_15 (pwire_11[15], swire_10[15], cwire_11[14], swire_11[14], cwire_11[15]);
fa f11_16 (pwire_11[16], swire_10[16], cwire_11[15], swire_11[15], cwire_11[16]);
fa f11_17 (pwire_11[17], swire_10[17], cwire_11[16], swire_11[16], cwire_11[17]);
fa f11_18 (pwire_11[18], swire_10[18], cwire_11[17], swire_11[17], cwire_11[18]);
fa f11_19 (pwire_11[19], swire_10[19], cwire_11[18], swire_11[18], cwire_11[19]);
fa f11_20 (pwire_11[20], swire_10[20], cwire_11[19], swire_11[19], cwire_11[20]);
fa f11_21 (pwire_11[21], swire_10[21], cwire_11[20], swire_11[20], cwire_11[21]);
fa f11_22 (pwire_11[22], swire_10[22], cwire_11[21], swire_11[21], cwire_11[22]);
fa f11_23 (pwire_11[23], swire_10[23], cwire_11[22], swire_11[22], cwire_11[23]);
fa f11_24 (pwire_11[24], swire_10[24], cwire_11[23], swire_11[23], cwire_11[24]);
fa f11_25 (pwire_11[25], swire_10[25], cwire_11[24], swire_11[24], cwire_11[25]);
fa f11_26 (pwire_11[26], swire_10[26], cwire_11[25], swire_11[25], cwire_11[26]);
fa f11_27 (pwire_11[27], swire_10[27], cwire_11[26], swire_11[26], cwire_11[27]);
fa f11_28 (pwire_11[28], swire_10[28], cwire_11[27], swire_11[27], cwire_11[28]);
fa f11_29 (pwire_11[29], swire_10[29], cwire_11[28], swire_11[28], cwire_11[29]);
fa f11_30 (pwire_11[30], swire_10[30], cwire_11[29], swire_11[29], cwire_11[30]);
fa f11_31 (pwire_11[31], swire_10[31], cwire_11[30], swire_11[30], cwire_11[31]);

//Stage11Padding
fa f11__1 (pwire_11[31], swire_10[32], cwire_11[31], swire_11[31], cwire_11[32]);
fa f11__2 (pwire_11[31], swire_10[33], cwire_11[32], swire_11[32], cwire_11[33]);
fa f11__3 (pwire_11[31], swire_10[34], cwire_11[33], swire_11[33], cwire_11[34]);
fa f11__4 (pwire_11[31], swire_10[35], cwire_11[34], swire_11[34], cwire_11[35]);
fa f11__5 (pwire_11[31], swire_10[36], cwire_11[35], swire_11[35], cwire_11[36]);
fa f11__6 (pwire_11[31], swire_10[37], cwire_11[36], swire_11[36], cwire_11[37]);
fa f11__7 (pwire_11[31], swire_10[38], cwire_11[37], swire_11[37], cwire_11[38]);
fa f11__8 (pwire_11[31], swire_10[39], cwire_11[38], swire_11[38], cwire_11[39]);
fa f11__9 (pwire_11[31], swire_10[40], cwire_11[39], swire_11[39], cwire_11[40]);
fa f11__10 (pwire_11[31], swire_10[41], cwire_11[40], swire_11[40], cwire_11[41]);
fa f11__11 (pwire_11[31], swire_10[42], cwire_11[41], swire_11[41], cwire_11[42]);
fa f11__12 (pwire_11[31], swire_10[43], cwire_11[42], swire_11[42], cwire_11[43]);
fa f11__13 (pwire_11[31], swire_10[44], cwire_11[43], swire_11[43], cwire_11[44]);
fa f11__14 (pwire_11[31], swire_10[45], cwire_11[44], swire_11[44], cwire_11[45]);
fa f11__15 (pwire_11[31], swire_10[46], cwire_11[45], swire_11[45], cwire_11[46]);
fa f11__16 (pwire_11[31], swire_10[47], cwire_11[46], swire_11[46], cwire_11[47]);
fa f11__17 (pwire_11[31], swire_10[48], cwire_11[47], swire_11[47], cwire_11[48]);
fa f11__18 (pwire_11[31], swire_10[49], cwire_11[48], swire_11[48], cwire_11[49]);
fa f11__19 (pwire_11[31], swire_10[50], cwire_11[49], swire_11[49], cwire_11[50]);
fa f11__20 (pwire_11[31], swire_10[51], cwire_11[50], swire_11[50], cwire_11[51]);
fa f11__21 (pwire_11[31], swire_10[52], cwire_11[51], swire_11[51], cwire_11[52]);

//Stage12 Partial Mul
ha f12(pwire_12[0], swire_11[0], mul[12], cwire_12[0]);
fa f12_1 (pwire_12[1], swire_11[1], cwire_12[0], swire_12[0], cwire_12[1]);
fa f12_2 (pwire_12[2], swire_11[2], cwire_12[1], swire_12[1], cwire_12[2]);
fa f12_3 (pwire_12[3], swire_11[3], cwire_12[2], swire_12[2], cwire_12[3]);
fa f12_4 (pwire_12[4], swire_11[4], cwire_12[3], swire_12[3], cwire_12[4]);
fa f12_5 (pwire_12[5], swire_11[5], cwire_12[4], swire_12[4], cwire_12[5]);
fa f12_6 (pwire_12[6], swire_11[6], cwire_12[5], swire_12[5], cwire_12[6]);
fa f12_7 (pwire_12[7], swire_11[7], cwire_12[6], swire_12[6], cwire_12[7]);
fa f12_8 (pwire_12[8], swire_11[8], cwire_12[7], swire_12[7], cwire_12[8]);
fa f12_9 (pwire_12[9], swire_11[9], cwire_12[8], swire_12[8], cwire_12[9]);
fa f12_10 (pwire_12[10], swire_11[10], cwire_12[9], swire_12[9], cwire_12[10]);
fa f12_11 (pwire_12[11], swire_11[11], cwire_12[10], swire_12[10], cwire_12[11]);
fa f12_12 (pwire_12[12], swire_11[12], cwire_12[11], swire_12[11], cwire_12[12]);
fa f12_13 (pwire_12[13], swire_11[13], cwire_12[12], swire_12[12], cwire_12[13]);
fa f12_14 (pwire_12[14], swire_11[14], cwire_12[13], swire_12[13], cwire_12[14]);
fa f12_15 (pwire_12[15], swire_11[15], cwire_12[14], swire_12[14], cwire_12[15]);
fa f12_16 (pwire_12[16], swire_11[16], cwire_12[15], swire_12[15], cwire_12[16]);
fa f12_17 (pwire_12[17], swire_11[17], cwire_12[16], swire_12[16], cwire_12[17]);
fa f12_18 (pwire_12[18], swire_11[18], cwire_12[17], swire_12[17], cwire_12[18]);
fa f12_19 (pwire_12[19], swire_11[19], cwire_12[18], swire_12[18], cwire_12[19]);
fa f12_20 (pwire_12[20], swire_11[20], cwire_12[19], swire_12[19], cwire_12[20]);
fa f12_21 (pwire_12[21], swire_11[21], cwire_12[20], swire_12[20], cwire_12[21]);
fa f12_22 (pwire_12[22], swire_11[22], cwire_12[21], swire_12[21], cwire_12[22]);
fa f12_23 (pwire_12[23], swire_11[23], cwire_12[22], swire_12[22], cwire_12[23]);
fa f12_24 (pwire_12[24], swire_11[24], cwire_12[23], swire_12[23], cwire_12[24]);
fa f12_25 (pwire_12[25], swire_11[25], cwire_12[24], swire_12[24], cwire_12[25]);
fa f12_26 (pwire_12[26], swire_11[26], cwire_12[25], swire_12[25], cwire_12[26]);
fa f12_27 (pwire_12[27], swire_11[27], cwire_12[26], swire_12[26], cwire_12[27]);
fa f12_28 (pwire_12[28], swire_11[28], cwire_12[27], swire_12[27], cwire_12[28]);
fa f12_29 (pwire_12[29], swire_11[29], cwire_12[28], swire_12[28], cwire_12[29]);
fa f12_30 (pwire_12[30], swire_11[30], cwire_12[29], swire_12[29], cwire_12[30]);
fa f12_31 (pwire_12[31], swire_11[31], cwire_12[30], swire_12[30], cwire_12[31]);

//Stage12Padding
fa f12__1 (pwire_12[31], swire_11[32], cwire_12[31], swire_12[31], cwire_12[32]);
fa f12__2 (pwire_12[31], swire_11[33], cwire_12[32], swire_12[32], cwire_12[33]);
fa f12__3 (pwire_12[31], swire_11[34], cwire_12[33], swire_12[33], cwire_12[34]);
fa f12__4 (pwire_12[31], swire_11[35], cwire_12[34], swire_12[34], cwire_12[35]);
fa f12__5 (pwire_12[31], swire_11[36], cwire_12[35], swire_12[35], cwire_12[36]);
fa f12__6 (pwire_12[31], swire_11[37], cwire_12[36], swire_12[36], cwire_12[37]);
fa f12__7 (pwire_12[31], swire_11[38], cwire_12[37], swire_12[37], cwire_12[38]);
fa f12__8 (pwire_12[31], swire_11[39], cwire_12[38], swire_12[38], cwire_12[39]);
fa f12__9 (pwire_12[31], swire_11[40], cwire_12[39], swire_12[39], cwire_12[40]);
fa f12__10 (pwire_12[31], swire_11[41], cwire_12[40], swire_12[40], cwire_12[41]);
fa f12__11 (pwire_12[31], swire_11[42], cwire_12[41], swire_12[41], cwire_12[42]);
fa f12__12 (pwire_12[31], swire_11[43], cwire_12[42], swire_12[42], cwire_12[43]);
fa f12__13 (pwire_12[31], swire_11[44], cwire_12[43], swire_12[43], cwire_12[44]);
fa f12__14 (pwire_12[31], swire_11[45], cwire_12[44], swire_12[44], cwire_12[45]);
fa f12__15 (pwire_12[31], swire_11[46], cwire_12[45], swire_12[45], cwire_12[46]);
fa f12__16 (pwire_12[31], swire_11[47], cwire_12[46], swire_12[46], cwire_12[47]);
fa f12__17 (pwire_12[31], swire_11[48], cwire_12[47], swire_12[47], cwire_12[48]);
fa f12__18 (pwire_12[31], swire_11[49], cwire_12[48], swire_12[48], cwire_12[49]);
fa f12__19 (pwire_12[31], swire_11[50], cwire_12[49], swire_12[49], cwire_12[50]);
fa f12__20 (pwire_12[31], swire_11[51], cwire_12[50], swire_12[50], cwire_12[51]);

//Stage13 Partial Mul
ha f13(pwire_13[0], swire_12[0], mul[13], cwire_13[0]);
fa f13_1 (pwire_13[1], swire_12[1], cwire_13[0], swire_13[0], cwire_13[1]);
fa f13_2 (pwire_13[2], swire_12[2], cwire_13[1], swire_13[1], cwire_13[2]);
fa f13_3 (pwire_13[3], swire_12[3], cwire_13[2], swire_13[2], cwire_13[3]);
fa f13_4 (pwire_13[4], swire_12[4], cwire_13[3], swire_13[3], cwire_13[4]);
fa f13_5 (pwire_13[5], swire_12[5], cwire_13[4], swire_13[4], cwire_13[5]);
fa f13_6 (pwire_13[6], swire_12[6], cwire_13[5], swire_13[5], cwire_13[6]);
fa f13_7 (pwire_13[7], swire_12[7], cwire_13[6], swire_13[6], cwire_13[7]);
fa f13_8 (pwire_13[8], swire_12[8], cwire_13[7], swire_13[7], cwire_13[8]);
fa f13_9 (pwire_13[9], swire_12[9], cwire_13[8], swire_13[8], cwire_13[9]);
fa f13_10 (pwire_13[10], swire_12[10], cwire_13[9], swire_13[9], cwire_13[10]);
fa f13_11 (pwire_13[11], swire_12[11], cwire_13[10], swire_13[10], cwire_13[11]);
fa f13_12 (pwire_13[12], swire_12[12], cwire_13[11], swire_13[11], cwire_13[12]);
fa f13_13 (pwire_13[13], swire_12[13], cwire_13[12], swire_13[12], cwire_13[13]);
fa f13_14 (pwire_13[14], swire_12[14], cwire_13[13], swire_13[13], cwire_13[14]);
fa f13_15 (pwire_13[15], swire_12[15], cwire_13[14], swire_13[14], cwire_13[15]);
fa f13_16 (pwire_13[16], swire_12[16], cwire_13[15], swire_13[15], cwire_13[16]);
fa f13_17 (pwire_13[17], swire_12[17], cwire_13[16], swire_13[16], cwire_13[17]);
fa f13_18 (pwire_13[18], swire_12[18], cwire_13[17], swire_13[17], cwire_13[18]);
fa f13_19 (pwire_13[19], swire_12[19], cwire_13[18], swire_13[18], cwire_13[19]);
fa f13_20 (pwire_13[20], swire_12[20], cwire_13[19], swire_13[19], cwire_13[20]);
fa f13_21 (pwire_13[21], swire_12[21], cwire_13[20], swire_13[20], cwire_13[21]);
fa f13_22 (pwire_13[22], swire_12[22], cwire_13[21], swire_13[21], cwire_13[22]);
fa f13_23 (pwire_13[23], swire_12[23], cwire_13[22], swire_13[22], cwire_13[23]);
fa f13_24 (pwire_13[24], swire_12[24], cwire_13[23], swire_13[23], cwire_13[24]);
fa f13_25 (pwire_13[25], swire_12[25], cwire_13[24], swire_13[24], cwire_13[25]);
fa f13_26 (pwire_13[26], swire_12[26], cwire_13[25], swire_13[25], cwire_13[26]);
fa f13_27 (pwire_13[27], swire_12[27], cwire_13[26], swire_13[26], cwire_13[27]);
fa f13_28 (pwire_13[28], swire_12[28], cwire_13[27], swire_13[27], cwire_13[28]);
fa f13_29 (pwire_13[29], swire_12[29], cwire_13[28], swire_13[28], cwire_13[29]);
fa f13_30 (pwire_13[30], swire_12[30], cwire_13[29], swire_13[29], cwire_13[30]);
fa f13_31 (pwire_13[31], swire_12[31], cwire_13[30], swire_13[30], cwire_13[31]);

//Stage13Padding
fa f13__1 (pwire_13[31], swire_12[32], cwire_13[31], swire_13[31], cwire_13[32]);
fa f13__2 (pwire_13[31], swire_12[33], cwire_13[32], swire_13[32], cwire_13[33]);
fa f13__3 (pwire_13[31], swire_12[34], cwire_13[33], swire_13[33], cwire_13[34]);
fa f13__4 (pwire_13[31], swire_12[35], cwire_13[34], swire_13[34], cwire_13[35]);
fa f13__5 (pwire_13[31], swire_12[36], cwire_13[35], swire_13[35], cwire_13[36]);
fa f13__6 (pwire_13[31], swire_12[37], cwire_13[36], swire_13[36], cwire_13[37]);
fa f13__7 (pwire_13[31], swire_12[38], cwire_13[37], swire_13[37], cwire_13[38]);
fa f13__8 (pwire_13[31], swire_12[39], cwire_13[38], swire_13[38], cwire_13[39]);
fa f13__9 (pwire_13[31], swire_12[40], cwire_13[39], swire_13[39], cwire_13[40]);
fa f13__10 (pwire_13[31], swire_12[41], cwire_13[40], swire_13[40], cwire_13[41]);
fa f13__11 (pwire_13[31], swire_12[42], cwire_13[41], swire_13[41], cwire_13[42]);
fa f13__12 (pwire_13[31], swire_12[43], cwire_13[42], swire_13[42], cwire_13[43]);
fa f13__13 (pwire_13[31], swire_12[44], cwire_13[43], swire_13[43], cwire_13[44]);
fa f13__14 (pwire_13[31], swire_12[45], cwire_13[44], swire_13[44], cwire_13[45]);
fa f13__15 (pwire_13[31], swire_12[46], cwire_13[45], swire_13[45], cwire_13[46]);
fa f13__16 (pwire_13[31], swire_12[47], cwire_13[46], swire_13[46], cwire_13[47]);
fa f13__17 (pwire_13[31], swire_12[48], cwire_13[47], swire_13[47], cwire_13[48]);
fa f13__18 (pwire_13[31], swire_12[49], cwire_13[48], swire_13[48], cwire_13[49]);
fa f13__19 (pwire_13[31], swire_12[50], cwire_13[49], swire_13[49], cwire_13[50]);

//Stage14 Partial Mul
ha f14(pwire_14[0], swire_13[0], mul[14], cwire_14[0]);
fa f14_1 (pwire_14[1], swire_13[1], cwire_14[0], swire_14[0], cwire_14[1]);
fa f14_2 (pwire_14[2], swire_13[2], cwire_14[1], swire_14[1], cwire_14[2]);
fa f14_3 (pwire_14[3], swire_13[3], cwire_14[2], swire_14[2], cwire_14[3]);
fa f14_4 (pwire_14[4], swire_13[4], cwire_14[3], swire_14[3], cwire_14[4]);
fa f14_5 (pwire_14[5], swire_13[5], cwire_14[4], swire_14[4], cwire_14[5]);
fa f14_6 (pwire_14[6], swire_13[6], cwire_14[5], swire_14[5], cwire_14[6]);
fa f14_7 (pwire_14[7], swire_13[7], cwire_14[6], swire_14[6], cwire_14[7]);
fa f14_8 (pwire_14[8], swire_13[8], cwire_14[7], swire_14[7], cwire_14[8]);
fa f14_9 (pwire_14[9], swire_13[9], cwire_14[8], swire_14[8], cwire_14[9]);
fa f14_10 (pwire_14[10], swire_13[10], cwire_14[9], swire_14[9], cwire_14[10]);
fa f14_11 (pwire_14[11], swire_13[11], cwire_14[10], swire_14[10], cwire_14[11]);
fa f14_12 (pwire_14[12], swire_13[12], cwire_14[11], swire_14[11], cwire_14[12]);
fa f14_13 (pwire_14[13], swire_13[13], cwire_14[12], swire_14[12], cwire_14[13]);
fa f14_14 (pwire_14[14], swire_13[14], cwire_14[13], swire_14[13], cwire_14[14]);
fa f14_15 (pwire_14[15], swire_13[15], cwire_14[14], swire_14[14], cwire_14[15]);
fa f14_16 (pwire_14[16], swire_13[16], cwire_14[15], swire_14[15], cwire_14[16]);
fa f14_17 (pwire_14[17], swire_13[17], cwire_14[16], swire_14[16], cwire_14[17]);
fa f14_18 (pwire_14[18], swire_13[18], cwire_14[17], swire_14[17], cwire_14[18]);
fa f14_19 (pwire_14[19], swire_13[19], cwire_14[18], swire_14[18], cwire_14[19]);
fa f14_20 (pwire_14[20], swire_13[20], cwire_14[19], swire_14[19], cwire_14[20]);
fa f14_21 (pwire_14[21], swire_13[21], cwire_14[20], swire_14[20], cwire_14[21]);
fa f14_22 (pwire_14[22], swire_13[22], cwire_14[21], swire_14[21], cwire_14[22]);
fa f14_23 (pwire_14[23], swire_13[23], cwire_14[22], swire_14[22], cwire_14[23]);
fa f14_24 (pwire_14[24], swire_13[24], cwire_14[23], swire_14[23], cwire_14[24]);
fa f14_25 (pwire_14[25], swire_13[25], cwire_14[24], swire_14[24], cwire_14[25]);
fa f14_26 (pwire_14[26], swire_13[26], cwire_14[25], swire_14[25], cwire_14[26]);
fa f14_27 (pwire_14[27], swire_13[27], cwire_14[26], swire_14[26], cwire_14[27]);
fa f14_28 (pwire_14[28], swire_13[28], cwire_14[27], swire_14[27], cwire_14[28]);
fa f14_29 (pwire_14[29], swire_13[29], cwire_14[28], swire_14[28], cwire_14[29]);
fa f14_30 (pwire_14[30], swire_13[30], cwire_14[29], swire_14[29], cwire_14[30]);
fa f14_31 (pwire_14[31], swire_13[31], cwire_14[30], swire_14[30], cwire_14[31]);

//Stage14Padding
fa f14__1 (pwire_14[31], swire_13[32], cwire_14[31], swire_14[31], cwire_14[32]);
fa f14__2 (pwire_14[31], swire_13[33], cwire_14[32], swire_14[32], cwire_14[33]);
fa f14__3 (pwire_14[31], swire_13[34], cwire_14[33], swire_14[33], cwire_14[34]);
fa f14__4 (pwire_14[31], swire_13[35], cwire_14[34], swire_14[34], cwire_14[35]);
fa f14__5 (pwire_14[31], swire_13[36], cwire_14[35], swire_14[35], cwire_14[36]);
fa f14__6 (pwire_14[31], swire_13[37], cwire_14[36], swire_14[36], cwire_14[37]);
fa f14__7 (pwire_14[31], swire_13[38], cwire_14[37], swire_14[37], cwire_14[38]);
fa f14__8 (pwire_14[31], swire_13[39], cwire_14[38], swire_14[38], cwire_14[39]);
fa f14__9 (pwire_14[31], swire_13[40], cwire_14[39], swire_14[39], cwire_14[40]);
fa f14__10 (pwire_14[31], swire_13[41], cwire_14[40], swire_14[40], cwire_14[41]);
fa f14__11 (pwire_14[31], swire_13[42], cwire_14[41], swire_14[41], cwire_14[42]);
fa f14__12 (pwire_14[31], swire_13[43], cwire_14[42], swire_14[42], cwire_14[43]);
fa f14__13 (pwire_14[31], swire_13[44], cwire_14[43], swire_14[43], cwire_14[44]);
fa f14__14 (pwire_14[31], swire_13[45], cwire_14[44], swire_14[44], cwire_14[45]);
fa f14__15 (pwire_14[31], swire_13[46], cwire_14[45], swire_14[45], cwire_14[46]);
fa f14__16 (pwire_14[31], swire_13[47], cwire_14[46], swire_14[46], cwire_14[47]);
fa f14__17 (pwire_14[31], swire_13[48], cwire_14[47], swire_14[47], cwire_14[48]);
fa f14__18 (pwire_14[31], swire_13[49], cwire_14[48], swire_14[48], cwire_14[49]);

//Stage15 Partial Mul
ha f15(pwire_15[0], swire_14[0], mul[15], cwire_15[0]);
fa f15_1 (pwire_15[1], swire_14[1], cwire_15[0], swire_15[0], cwire_15[1]);
fa f15_2 (pwire_15[2], swire_14[2], cwire_15[1], swire_15[1], cwire_15[2]);
fa f15_3 (pwire_15[3], swire_14[3], cwire_15[2], swire_15[2], cwire_15[3]);
fa f15_4 (pwire_15[4], swire_14[4], cwire_15[3], swire_15[3], cwire_15[4]);
fa f15_5 (pwire_15[5], swire_14[5], cwire_15[4], swire_15[4], cwire_15[5]);
fa f15_6 (pwire_15[6], swire_14[6], cwire_15[5], swire_15[5], cwire_15[6]);
fa f15_7 (pwire_15[7], swire_14[7], cwire_15[6], swire_15[6], cwire_15[7]);
fa f15_8 (pwire_15[8], swire_14[8], cwire_15[7], swire_15[7], cwire_15[8]);
fa f15_9 (pwire_15[9], swire_14[9], cwire_15[8], swire_15[8], cwire_15[9]);
fa f15_10 (pwire_15[10], swire_14[10], cwire_15[9], swire_15[9], cwire_15[10]);
fa f15_11 (pwire_15[11], swire_14[11], cwire_15[10], swire_15[10], cwire_15[11]);
fa f15_12 (pwire_15[12], swire_14[12], cwire_15[11], swire_15[11], cwire_15[12]);
fa f15_13 (pwire_15[13], swire_14[13], cwire_15[12], swire_15[12], cwire_15[13]);
fa f15_14 (pwire_15[14], swire_14[14], cwire_15[13], swire_15[13], cwire_15[14]);
fa f15_15 (pwire_15[15], swire_14[15], cwire_15[14], swire_15[14], cwire_15[15]);
fa f15_16 (pwire_15[16], swire_14[16], cwire_15[15], swire_15[15], cwire_15[16]);
fa f15_17 (pwire_15[17], swire_14[17], cwire_15[16], swire_15[16], cwire_15[17]);
fa f15_18 (pwire_15[18], swire_14[18], cwire_15[17], swire_15[17], cwire_15[18]);
fa f15_19 (pwire_15[19], swire_14[19], cwire_15[18], swire_15[18], cwire_15[19]);
fa f15_20 (pwire_15[20], swire_14[20], cwire_15[19], swire_15[19], cwire_15[20]);
fa f15_21 (pwire_15[21], swire_14[21], cwire_15[20], swire_15[20], cwire_15[21]);
fa f15_22 (pwire_15[22], swire_14[22], cwire_15[21], swire_15[21], cwire_15[22]);
fa f15_23 (pwire_15[23], swire_14[23], cwire_15[22], swire_15[22], cwire_15[23]);
fa f15_24 (pwire_15[24], swire_14[24], cwire_15[23], swire_15[23], cwire_15[24]);
fa f15_25 (pwire_15[25], swire_14[25], cwire_15[24], swire_15[24], cwire_15[25]);
fa f15_26 (pwire_15[26], swire_14[26], cwire_15[25], swire_15[25], cwire_15[26]);
fa f15_27 (pwire_15[27], swire_14[27], cwire_15[26], swire_15[26], cwire_15[27]);
fa f15_28 (pwire_15[28], swire_14[28], cwire_15[27], swire_15[27], cwire_15[28]);
fa f15_29 (pwire_15[29], swire_14[29], cwire_15[28], swire_15[28], cwire_15[29]);
fa f15_30 (pwire_15[30], swire_14[30], cwire_15[29], swire_15[29], cwire_15[30]);
fa f15_31 (pwire_15[31], swire_14[31], cwire_15[30], swire_15[30], cwire_15[31]);

//Stage15Padding
fa f15__1 (pwire_15[31], swire_14[32], cwire_15[31], swire_15[31], cwire_15[32]);
fa f15__2 (pwire_15[31], swire_14[33], cwire_15[32], swire_15[32], cwire_15[33]);
fa f15__3 (pwire_15[31], swire_14[34], cwire_15[33], swire_15[33], cwire_15[34]);
fa f15__4 (pwire_15[31], swire_14[35], cwire_15[34], swire_15[34], cwire_15[35]);
fa f15__5 (pwire_15[31], swire_14[36], cwire_15[35], swire_15[35], cwire_15[36]);
fa f15__6 (pwire_15[31], swire_14[37], cwire_15[36], swire_15[36], cwire_15[37]);
fa f15__7 (pwire_15[31], swire_14[38], cwire_15[37], swire_15[37], cwire_15[38]);
fa f15__8 (pwire_15[31], swire_14[39], cwire_15[38], swire_15[38], cwire_15[39]);
fa f15__9 (pwire_15[31], swire_14[40], cwire_15[39], swire_15[39], cwire_15[40]);
fa f15__10 (pwire_15[31], swire_14[41], cwire_15[40], swire_15[40], cwire_15[41]);
fa f15__11 (pwire_15[31], swire_14[42], cwire_15[41], swire_15[41], cwire_15[42]);
fa f15__12 (pwire_15[31], swire_14[43], cwire_15[42], swire_15[42], cwire_15[43]);
fa f15__13 (pwire_15[31], swire_14[44], cwire_15[43], swire_15[43], cwire_15[44]);
fa f15__14 (pwire_15[31], swire_14[45], cwire_15[44], swire_15[44], cwire_15[45]);
fa f15__15 (pwire_15[31], swire_14[46], cwire_15[45], swire_15[45], cwire_15[46]);
fa f15__16 (pwire_15[31], swire_14[47], cwire_15[46], swire_15[46], cwire_15[47]);
fa f15__17 (pwire_15[31], swire_14[48], cwire_15[47], swire_15[47], cwire_15[48]);

//Stage16 Partial Mul
ha f16(pwire_16[0], swire_15[0], mul[16], cwire_16[0]);
fa f16_1 (pwire_16[1], swire_15[1], cwire_16[0], swire_16[0], cwire_16[1]);
fa f16_2 (pwire_16[2], swire_15[2], cwire_16[1], swire_16[1], cwire_16[2]);
fa f16_3 (pwire_16[3], swire_15[3], cwire_16[2], swire_16[2], cwire_16[3]);
fa f16_4 (pwire_16[4], swire_15[4], cwire_16[3], swire_16[3], cwire_16[4]);
fa f16_5 (pwire_16[5], swire_15[5], cwire_16[4], swire_16[4], cwire_16[5]);
fa f16_6 (pwire_16[6], swire_15[6], cwire_16[5], swire_16[5], cwire_16[6]);
fa f16_7 (pwire_16[7], swire_15[7], cwire_16[6], swire_16[6], cwire_16[7]);
fa f16_8 (pwire_16[8], swire_15[8], cwire_16[7], swire_16[7], cwire_16[8]);
fa f16_9 (pwire_16[9], swire_15[9], cwire_16[8], swire_16[8], cwire_16[9]);
fa f16_10 (pwire_16[10], swire_15[10], cwire_16[9], swire_16[9], cwire_16[10]);
fa f16_11 (pwire_16[11], swire_15[11], cwire_16[10], swire_16[10], cwire_16[11]);
fa f16_12 (pwire_16[12], swire_15[12], cwire_16[11], swire_16[11], cwire_16[12]);
fa f16_13 (pwire_16[13], swire_15[13], cwire_16[12], swire_16[12], cwire_16[13]);
fa f16_14 (pwire_16[14], swire_15[14], cwire_16[13], swire_16[13], cwire_16[14]);
fa f16_15 (pwire_16[15], swire_15[15], cwire_16[14], swire_16[14], cwire_16[15]);
fa f16_16 (pwire_16[16], swire_15[16], cwire_16[15], swire_16[15], cwire_16[16]);
fa f16_17 (pwire_16[17], swire_15[17], cwire_16[16], swire_16[16], cwire_16[17]);
fa f16_18 (pwire_16[18], swire_15[18], cwire_16[17], swire_16[17], cwire_16[18]);
fa f16_19 (pwire_16[19], swire_15[19], cwire_16[18], swire_16[18], cwire_16[19]);
fa f16_20 (pwire_16[20], swire_15[20], cwire_16[19], swire_16[19], cwire_16[20]);
fa f16_21 (pwire_16[21], swire_15[21], cwire_16[20], swire_16[20], cwire_16[21]);
fa f16_22 (pwire_16[22], swire_15[22], cwire_16[21], swire_16[21], cwire_16[22]);
fa f16_23 (pwire_16[23], swire_15[23], cwire_16[22], swire_16[22], cwire_16[23]);
fa f16_24 (pwire_16[24], swire_15[24], cwire_16[23], swire_16[23], cwire_16[24]);
fa f16_25 (pwire_16[25], swire_15[25], cwire_16[24], swire_16[24], cwire_16[25]);
fa f16_26 (pwire_16[26], swire_15[26], cwire_16[25], swire_16[25], cwire_16[26]);
fa f16_27 (pwire_16[27], swire_15[27], cwire_16[26], swire_16[26], cwire_16[27]);
fa f16_28 (pwire_16[28], swire_15[28], cwire_16[27], swire_16[27], cwire_16[28]);
fa f16_29 (pwire_16[29], swire_15[29], cwire_16[28], swire_16[28], cwire_16[29]);
fa f16_30 (pwire_16[30], swire_15[30], cwire_16[29], swire_16[29], cwire_16[30]);
fa f16_31 (pwire_16[31], swire_15[31], cwire_16[30], swire_16[30], cwire_16[31]);

//Stage16Padding
fa f16__1 (pwire_16[31], swire_15[32], cwire_16[31], swire_16[31], cwire_16[32]);
fa f16__2 (pwire_16[31], swire_15[33], cwire_16[32], swire_16[32], cwire_16[33]);
fa f16__3 (pwire_16[31], swire_15[34], cwire_16[33], swire_16[33], cwire_16[34]);
fa f16__4 (pwire_16[31], swire_15[35], cwire_16[34], swire_16[34], cwire_16[35]);
fa f16__5 (pwire_16[31], swire_15[36], cwire_16[35], swire_16[35], cwire_16[36]);
fa f16__6 (pwire_16[31], swire_15[37], cwire_16[36], swire_16[36], cwire_16[37]);
fa f16__7 (pwire_16[31], swire_15[38], cwire_16[37], swire_16[37], cwire_16[38]);
fa f16__8 (pwire_16[31], swire_15[39], cwire_16[38], swire_16[38], cwire_16[39]);
fa f16__9 (pwire_16[31], swire_15[40], cwire_16[39], swire_16[39], cwire_16[40]);
fa f16__10 (pwire_16[31], swire_15[41], cwire_16[40], swire_16[40], cwire_16[41]);
fa f16__11 (pwire_16[31], swire_15[42], cwire_16[41], swire_16[41], cwire_16[42]);
fa f16__12 (pwire_16[31], swire_15[43], cwire_16[42], swire_16[42], cwire_16[43]);
fa f16__13 (pwire_16[31], swire_15[44], cwire_16[43], swire_16[43], cwire_16[44]);
fa f16__14 (pwire_16[31], swire_15[45], cwire_16[44], swire_16[44], cwire_16[45]);
fa f16__15 (pwire_16[31], swire_15[46], cwire_16[45], swire_16[45], cwire_16[46]);
fa f16__16 (pwire_16[31], swire_15[47], cwire_16[46], swire_16[46], cwire_16[47]);

//Stage17 Partial Mul
ha f17(pwire_17[0], swire_16[0], mul[17], cwire_17[0]);
fa f17_1 (pwire_17[1], swire_16[1], cwire_17[0], swire_17[0], cwire_17[1]);
fa f17_2 (pwire_17[2], swire_16[2], cwire_17[1], swire_17[1], cwire_17[2]);
fa f17_3 (pwire_17[3], swire_16[3], cwire_17[2], swire_17[2], cwire_17[3]);
fa f17_4 (pwire_17[4], swire_16[4], cwire_17[3], swire_17[3], cwire_17[4]);
fa f17_5 (pwire_17[5], swire_16[5], cwire_17[4], swire_17[4], cwire_17[5]);
fa f17_6 (pwire_17[6], swire_16[6], cwire_17[5], swire_17[5], cwire_17[6]);
fa f17_7 (pwire_17[7], swire_16[7], cwire_17[6], swire_17[6], cwire_17[7]);
fa f17_8 (pwire_17[8], swire_16[8], cwire_17[7], swire_17[7], cwire_17[8]);
fa f17_9 (pwire_17[9], swire_16[9], cwire_17[8], swire_17[8], cwire_17[9]);
fa f17_10 (pwire_17[10], swire_16[10], cwire_17[9], swire_17[9], cwire_17[10]);
fa f17_11 (pwire_17[11], swire_16[11], cwire_17[10], swire_17[10], cwire_17[11]);
fa f17_12 (pwire_17[12], swire_16[12], cwire_17[11], swire_17[11], cwire_17[12]);
fa f17_13 (pwire_17[13], swire_16[13], cwire_17[12], swire_17[12], cwire_17[13]);
fa f17_14 (pwire_17[14], swire_16[14], cwire_17[13], swire_17[13], cwire_17[14]);
fa f17_15 (pwire_17[15], swire_16[15], cwire_17[14], swire_17[14], cwire_17[15]);
fa f17_16 (pwire_17[16], swire_16[16], cwire_17[15], swire_17[15], cwire_17[16]);
fa f17_17 (pwire_17[17], swire_16[17], cwire_17[16], swire_17[16], cwire_17[17]);
fa f17_18 (pwire_17[18], swire_16[18], cwire_17[17], swire_17[17], cwire_17[18]);
fa f17_19 (pwire_17[19], swire_16[19], cwire_17[18], swire_17[18], cwire_17[19]);
fa f17_20 (pwire_17[20], swire_16[20], cwire_17[19], swire_17[19], cwire_17[20]);
fa f17_21 (pwire_17[21], swire_16[21], cwire_17[20], swire_17[20], cwire_17[21]);
fa f17_22 (pwire_17[22], swire_16[22], cwire_17[21], swire_17[21], cwire_17[22]);
fa f17_23 (pwire_17[23], swire_16[23], cwire_17[22], swire_17[22], cwire_17[23]);
fa f17_24 (pwire_17[24], swire_16[24], cwire_17[23], swire_17[23], cwire_17[24]);
fa f17_25 (pwire_17[25], swire_16[25], cwire_17[24], swire_17[24], cwire_17[25]);
fa f17_26 (pwire_17[26], swire_16[26], cwire_17[25], swire_17[25], cwire_17[26]);
fa f17_27 (pwire_17[27], swire_16[27], cwire_17[26], swire_17[26], cwire_17[27]);
fa f17_28 (pwire_17[28], swire_16[28], cwire_17[27], swire_17[27], cwire_17[28]);
fa f17_29 (pwire_17[29], swire_16[29], cwire_17[28], swire_17[28], cwire_17[29]);
fa f17_30 (pwire_17[30], swire_16[30], cwire_17[29], swire_17[29], cwire_17[30]);
fa f17_31 (pwire_17[31], swire_16[31], cwire_17[30], swire_17[30], cwire_17[31]);

//Stage17Padding
fa f17__1 (pwire_17[31], swire_16[32], cwire_17[31], swire_17[31], cwire_17[32]);
fa f17__2 (pwire_17[31], swire_16[33], cwire_17[32], swire_17[32], cwire_17[33]);
fa f17__3 (pwire_17[31], swire_16[34], cwire_17[33], swire_17[33], cwire_17[34]);
fa f17__4 (pwire_17[31], swire_16[35], cwire_17[34], swire_17[34], cwire_17[35]);
fa f17__5 (pwire_17[31], swire_16[36], cwire_17[35], swire_17[35], cwire_17[36]);
fa f17__6 (pwire_17[31], swire_16[37], cwire_17[36], swire_17[36], cwire_17[37]);
fa f17__7 (pwire_17[31], swire_16[38], cwire_17[37], swire_17[37], cwire_17[38]);
fa f17__8 (pwire_17[31], swire_16[39], cwire_17[38], swire_17[38], cwire_17[39]);
fa f17__9 (pwire_17[31], swire_16[40], cwire_17[39], swire_17[39], cwire_17[40]);
fa f17__10 (pwire_17[31], swire_16[41], cwire_17[40], swire_17[40], cwire_17[41]);
fa f17__11 (pwire_17[31], swire_16[42], cwire_17[41], swire_17[41], cwire_17[42]);
fa f17__12 (pwire_17[31], swire_16[43], cwire_17[42], swire_17[42], cwire_17[43]);
fa f17__13 (pwire_17[31], swire_16[44], cwire_17[43], swire_17[43], cwire_17[44]);
fa f17__14 (pwire_17[31], swire_16[45], cwire_17[44], swire_17[44], cwire_17[45]);
fa f17__15 (pwire_17[31], swire_16[46], cwire_17[45], swire_17[45], cwire_17[46]);

//Stage18 Partial Mul
ha f18(pwire_18[0], swire_17[0], mul[18], cwire_18[0]);
fa f18_1 (pwire_18[1], swire_17[1], cwire_18[0], swire_18[0], cwire_18[1]);
fa f18_2 (pwire_18[2], swire_17[2], cwire_18[1], swire_18[1], cwire_18[2]);
fa f18_3 (pwire_18[3], swire_17[3], cwire_18[2], swire_18[2], cwire_18[3]);
fa f18_4 (pwire_18[4], swire_17[4], cwire_18[3], swire_18[3], cwire_18[4]);
fa f18_5 (pwire_18[5], swire_17[5], cwire_18[4], swire_18[4], cwire_18[5]);
fa f18_6 (pwire_18[6], swire_17[6], cwire_18[5], swire_18[5], cwire_18[6]);
fa f18_7 (pwire_18[7], swire_17[7], cwire_18[6], swire_18[6], cwire_18[7]);
fa f18_8 (pwire_18[8], swire_17[8], cwire_18[7], swire_18[7], cwire_18[8]);
fa f18_9 (pwire_18[9], swire_17[9], cwire_18[8], swire_18[8], cwire_18[9]);
fa f18_10 (pwire_18[10], swire_17[10], cwire_18[9], swire_18[9], cwire_18[10]);
fa f18_11 (pwire_18[11], swire_17[11], cwire_18[10], swire_18[10], cwire_18[11]);
fa f18_12 (pwire_18[12], swire_17[12], cwire_18[11], swire_18[11], cwire_18[12]);
fa f18_13 (pwire_18[13], swire_17[13], cwire_18[12], swire_18[12], cwire_18[13]);
fa f18_14 (pwire_18[14], swire_17[14], cwire_18[13], swire_18[13], cwire_18[14]);
fa f18_15 (pwire_18[15], swire_17[15], cwire_18[14], swire_18[14], cwire_18[15]);
fa f18_16 (pwire_18[16], swire_17[16], cwire_18[15], swire_18[15], cwire_18[16]);
fa f18_17 (pwire_18[17], swire_17[17], cwire_18[16], swire_18[16], cwire_18[17]);
fa f18_18 (pwire_18[18], swire_17[18], cwire_18[17], swire_18[17], cwire_18[18]);
fa f18_19 (pwire_18[19], swire_17[19], cwire_18[18], swire_18[18], cwire_18[19]);
fa f18_20 (pwire_18[20], swire_17[20], cwire_18[19], swire_18[19], cwire_18[20]);
fa f18_21 (pwire_18[21], swire_17[21], cwire_18[20], swire_18[20], cwire_18[21]);
fa f18_22 (pwire_18[22], swire_17[22], cwire_18[21], swire_18[21], cwire_18[22]);
fa f18_23 (pwire_18[23], swire_17[23], cwire_18[22], swire_18[22], cwire_18[23]);
fa f18_24 (pwire_18[24], swire_17[24], cwire_18[23], swire_18[23], cwire_18[24]);
fa f18_25 (pwire_18[25], swire_17[25], cwire_18[24], swire_18[24], cwire_18[25]);
fa f18_26 (pwire_18[26], swire_17[26], cwire_18[25], swire_18[25], cwire_18[26]);
fa f18_27 (pwire_18[27], swire_17[27], cwire_18[26], swire_18[26], cwire_18[27]);
fa f18_28 (pwire_18[28], swire_17[28], cwire_18[27], swire_18[27], cwire_18[28]);
fa f18_29 (pwire_18[29], swire_17[29], cwire_18[28], swire_18[28], cwire_18[29]);
fa f18_30 (pwire_18[30], swire_17[30], cwire_18[29], swire_18[29], cwire_18[30]);
fa f18_31 (pwire_18[31], swire_17[31], cwire_18[30], swire_18[30], cwire_18[31]);

//Stage18Padding
fa f18__1 (pwire_18[31], swire_17[32], cwire_18[31], swire_18[31], cwire_18[32]);
fa f18__2 (pwire_18[31], swire_17[33], cwire_18[32], swire_18[32], cwire_18[33]);
fa f18__3 (pwire_18[31], swire_17[34], cwire_18[33], swire_18[33], cwire_18[34]);
fa f18__4 (pwire_18[31], swire_17[35], cwire_18[34], swire_18[34], cwire_18[35]);
fa f18__5 (pwire_18[31], swire_17[36], cwire_18[35], swire_18[35], cwire_18[36]);
fa f18__6 (pwire_18[31], swire_17[37], cwire_18[36], swire_18[36], cwire_18[37]);
fa f18__7 (pwire_18[31], swire_17[38], cwire_18[37], swire_18[37], cwire_18[38]);
fa f18__8 (pwire_18[31], swire_17[39], cwire_18[38], swire_18[38], cwire_18[39]);
fa f18__9 (pwire_18[31], swire_17[40], cwire_18[39], swire_18[39], cwire_18[40]);
fa f18__10 (pwire_18[31], swire_17[41], cwire_18[40], swire_18[40], cwire_18[41]);
fa f18__11 (pwire_18[31], swire_17[42], cwire_18[41], swire_18[41], cwire_18[42]);
fa f18__12 (pwire_18[31], swire_17[43], cwire_18[42], swire_18[42], cwire_18[43]);
fa f18__13 (pwire_18[31], swire_17[44], cwire_18[43], swire_18[43], cwire_18[44]);
fa f18__14 (pwire_18[31], swire_17[45], cwire_18[44], swire_18[44], cwire_18[45]);

//Stage19 Partial Mul
ha f19(pwire_19[0], swire_18[0], mul[19], cwire_19[0]);
fa f19_1 (pwire_19[1], swire_18[1], cwire_19[0], swire_19[0], cwire_19[1]);
fa f19_2 (pwire_19[2], swire_18[2], cwire_19[1], swire_19[1], cwire_19[2]);
fa f19_3 (pwire_19[3], swire_18[3], cwire_19[2], swire_19[2], cwire_19[3]);
fa f19_4 (pwire_19[4], swire_18[4], cwire_19[3], swire_19[3], cwire_19[4]);
fa f19_5 (pwire_19[5], swire_18[5], cwire_19[4], swire_19[4], cwire_19[5]);
fa f19_6 (pwire_19[6], swire_18[6], cwire_19[5], swire_19[5], cwire_19[6]);
fa f19_7 (pwire_19[7], swire_18[7], cwire_19[6], swire_19[6], cwire_19[7]);
fa f19_8 (pwire_19[8], swire_18[8], cwire_19[7], swire_19[7], cwire_19[8]);
fa f19_9 (pwire_19[9], swire_18[9], cwire_19[8], swire_19[8], cwire_19[9]);
fa f19_10 (pwire_19[10], swire_18[10], cwire_19[9], swire_19[9], cwire_19[10]);
fa f19_11 (pwire_19[11], swire_18[11], cwire_19[10], swire_19[10], cwire_19[11]);
fa f19_12 (pwire_19[12], swire_18[12], cwire_19[11], swire_19[11], cwire_19[12]);
fa f19_13 (pwire_19[13], swire_18[13], cwire_19[12], swire_19[12], cwire_19[13]);
fa f19_14 (pwire_19[14], swire_18[14], cwire_19[13], swire_19[13], cwire_19[14]);
fa f19_15 (pwire_19[15], swire_18[15], cwire_19[14], swire_19[14], cwire_19[15]);
fa f19_16 (pwire_19[16], swire_18[16], cwire_19[15], swire_19[15], cwire_19[16]);
fa f19_17 (pwire_19[17], swire_18[17], cwire_19[16], swire_19[16], cwire_19[17]);
fa f19_18 (pwire_19[18], swire_18[18], cwire_19[17], swire_19[17], cwire_19[18]);
fa f19_19 (pwire_19[19], swire_18[19], cwire_19[18], swire_19[18], cwire_19[19]);
fa f19_20 (pwire_19[20], swire_18[20], cwire_19[19], swire_19[19], cwire_19[20]);
fa f19_21 (pwire_19[21], swire_18[21], cwire_19[20], swire_19[20], cwire_19[21]);
fa f19_22 (pwire_19[22], swire_18[22], cwire_19[21], swire_19[21], cwire_19[22]);
fa f19_23 (pwire_19[23], swire_18[23], cwire_19[22], swire_19[22], cwire_19[23]);
fa f19_24 (pwire_19[24], swire_18[24], cwire_19[23], swire_19[23], cwire_19[24]);
fa f19_25 (pwire_19[25], swire_18[25], cwire_19[24], swire_19[24], cwire_19[25]);
fa f19_26 (pwire_19[26], swire_18[26], cwire_19[25], swire_19[25], cwire_19[26]);
fa f19_27 (pwire_19[27], swire_18[27], cwire_19[26], swire_19[26], cwire_19[27]);
fa f19_28 (pwire_19[28], swire_18[28], cwire_19[27], swire_19[27], cwire_19[28]);
fa f19_29 (pwire_19[29], swire_18[29], cwire_19[28], swire_19[28], cwire_19[29]);
fa f19_30 (pwire_19[30], swire_18[30], cwire_19[29], swire_19[29], cwire_19[30]);
fa f19_31 (pwire_19[31], swire_18[31], cwire_19[30], swire_19[30], cwire_19[31]);

//Stage19Padding
fa f19__1 (pwire_19[31], swire_18[32], cwire_19[31], swire_19[31], cwire_19[32]);
fa f19__2 (pwire_19[31], swire_18[33], cwire_19[32], swire_19[32], cwire_19[33]);
fa f19__3 (pwire_19[31], swire_18[34], cwire_19[33], swire_19[33], cwire_19[34]);
fa f19__4 (pwire_19[31], swire_18[35], cwire_19[34], swire_19[34], cwire_19[35]);
fa f19__5 (pwire_19[31], swire_18[36], cwire_19[35], swire_19[35], cwire_19[36]);
fa f19__6 (pwire_19[31], swire_18[37], cwire_19[36], swire_19[36], cwire_19[37]);
fa f19__7 (pwire_19[31], swire_18[38], cwire_19[37], swire_19[37], cwire_19[38]);
fa f19__8 (pwire_19[31], swire_18[39], cwire_19[38], swire_19[38], cwire_19[39]);
fa f19__9 (pwire_19[31], swire_18[40], cwire_19[39], swire_19[39], cwire_19[40]);
fa f19__10 (pwire_19[31], swire_18[41], cwire_19[40], swire_19[40], cwire_19[41]);
fa f19__11 (pwire_19[31], swire_18[42], cwire_19[41], swire_19[41], cwire_19[42]);
fa f19__12 (pwire_19[31], swire_18[43], cwire_19[42], swire_19[42], cwire_19[43]);
fa f19__13 (pwire_19[31], swire_18[44], cwire_19[43], swire_19[43], cwire_19[44]);

//Stage20 Partial Mul
ha f20(pwire_20[0], swire_19[0], mul[20], cwire_20[0]);
fa f20_1 (pwire_20[1], swire_19[1], cwire_20[0], swire_20[0], cwire_20[1]);
fa f20_2 (pwire_20[2], swire_19[2], cwire_20[1], swire_20[1], cwire_20[2]);
fa f20_3 (pwire_20[3], swire_19[3], cwire_20[2], swire_20[2], cwire_20[3]);
fa f20_4 (pwire_20[4], swire_19[4], cwire_20[3], swire_20[3], cwire_20[4]);
fa f20_5 (pwire_20[5], swire_19[5], cwire_20[4], swire_20[4], cwire_20[5]);
fa f20_6 (pwire_20[6], swire_19[6], cwire_20[5], swire_20[5], cwire_20[6]);
fa f20_7 (pwire_20[7], swire_19[7], cwire_20[6], swire_20[6], cwire_20[7]);
fa f20_8 (pwire_20[8], swire_19[8], cwire_20[7], swire_20[7], cwire_20[8]);
fa f20_9 (pwire_20[9], swire_19[9], cwire_20[8], swire_20[8], cwire_20[9]);
fa f20_10 (pwire_20[10], swire_19[10], cwire_20[9], swire_20[9], cwire_20[10]);
fa f20_11 (pwire_20[11], swire_19[11], cwire_20[10], swire_20[10], cwire_20[11]);
fa f20_12 (pwire_20[12], swire_19[12], cwire_20[11], swire_20[11], cwire_20[12]);
fa f20_13 (pwire_20[13], swire_19[13], cwire_20[12], swire_20[12], cwire_20[13]);
fa f20_14 (pwire_20[14], swire_19[14], cwire_20[13], swire_20[13], cwire_20[14]);
fa f20_15 (pwire_20[15], swire_19[15], cwire_20[14], swire_20[14], cwire_20[15]);
fa f20_16 (pwire_20[16], swire_19[16], cwire_20[15], swire_20[15], cwire_20[16]);
fa f20_17 (pwire_20[17], swire_19[17], cwire_20[16], swire_20[16], cwire_20[17]);
fa f20_18 (pwire_20[18], swire_19[18], cwire_20[17], swire_20[17], cwire_20[18]);
fa f20_19 (pwire_20[19], swire_19[19], cwire_20[18], swire_20[18], cwire_20[19]);
fa f20_20 (pwire_20[20], swire_19[20], cwire_20[19], swire_20[19], cwire_20[20]);
fa f20_21 (pwire_20[21], swire_19[21], cwire_20[20], swire_20[20], cwire_20[21]);
fa f20_22 (pwire_20[22], swire_19[22], cwire_20[21], swire_20[21], cwire_20[22]);
fa f20_23 (pwire_20[23], swire_19[23], cwire_20[22], swire_20[22], cwire_20[23]);
fa f20_24 (pwire_20[24], swire_19[24], cwire_20[23], swire_20[23], cwire_20[24]);
fa f20_25 (pwire_20[25], swire_19[25], cwire_20[24], swire_20[24], cwire_20[25]);
fa f20_26 (pwire_20[26], swire_19[26], cwire_20[25], swire_20[25], cwire_20[26]);
fa f20_27 (pwire_20[27], swire_19[27], cwire_20[26], swire_20[26], cwire_20[27]);
fa f20_28 (pwire_20[28], swire_19[28], cwire_20[27], swire_20[27], cwire_20[28]);
fa f20_29 (pwire_20[29], swire_19[29], cwire_20[28], swire_20[28], cwire_20[29]);
fa f20_30 (pwire_20[30], swire_19[30], cwire_20[29], swire_20[29], cwire_20[30]);
fa f20_31 (pwire_20[31], swire_19[31], cwire_20[30], swire_20[30], cwire_20[31]);

//Stage20Padding
fa f20__1 (pwire_20[31], swire_19[32], cwire_20[31], swire_20[31], cwire_20[32]);
fa f20__2 (pwire_20[31], swire_19[33], cwire_20[32], swire_20[32], cwire_20[33]);
fa f20__3 (pwire_20[31], swire_19[34], cwire_20[33], swire_20[33], cwire_20[34]);
fa f20__4 (pwire_20[31], swire_19[35], cwire_20[34], swire_20[34], cwire_20[35]);
fa f20__5 (pwire_20[31], swire_19[36], cwire_20[35], swire_20[35], cwire_20[36]);
fa f20__6 (pwire_20[31], swire_19[37], cwire_20[36], swire_20[36], cwire_20[37]);
fa f20__7 (pwire_20[31], swire_19[38], cwire_20[37], swire_20[37], cwire_20[38]);
fa f20__8 (pwire_20[31], swire_19[39], cwire_20[38], swire_20[38], cwire_20[39]);
fa f20__9 (pwire_20[31], swire_19[40], cwire_20[39], swire_20[39], cwire_20[40]);
fa f20__10 (pwire_20[31], swire_19[41], cwire_20[40], swire_20[40], cwire_20[41]);
fa f20__11 (pwire_20[31], swire_19[42], cwire_20[41], swire_20[41], cwire_20[42]);
fa f20__12 (pwire_20[31], swire_19[43], cwire_20[42], swire_20[42], cwire_20[43]);

//Stage21 Partial Mul
ha f21(pwire_21[0], swire_20[0], mul[21], cwire_21[0]);
fa f21_1 (pwire_21[1], swire_20[1], cwire_21[0], swire_21[0], cwire_21[1]);
fa f21_2 (pwire_21[2], swire_20[2], cwire_21[1], swire_21[1], cwire_21[2]);
fa f21_3 (pwire_21[3], swire_20[3], cwire_21[2], swire_21[2], cwire_21[3]);
fa f21_4 (pwire_21[4], swire_20[4], cwire_21[3], swire_21[3], cwire_21[4]);
fa f21_5 (pwire_21[5], swire_20[5], cwire_21[4], swire_21[4], cwire_21[5]);
fa f21_6 (pwire_21[6], swire_20[6], cwire_21[5], swire_21[5], cwire_21[6]);
fa f21_7 (pwire_21[7], swire_20[7], cwire_21[6], swire_21[6], cwire_21[7]);
fa f21_8 (pwire_21[8], swire_20[8], cwire_21[7], swire_21[7], cwire_21[8]);
fa f21_9 (pwire_21[9], swire_20[9], cwire_21[8], swire_21[8], cwire_21[9]);
fa f21_10 (pwire_21[10], swire_20[10], cwire_21[9], swire_21[9], cwire_21[10]);
fa f21_11 (pwire_21[11], swire_20[11], cwire_21[10], swire_21[10], cwire_21[11]);
fa f21_12 (pwire_21[12], swire_20[12], cwire_21[11], swire_21[11], cwire_21[12]);
fa f21_13 (pwire_21[13], swire_20[13], cwire_21[12], swire_21[12], cwire_21[13]);
fa f21_14 (pwire_21[14], swire_20[14], cwire_21[13], swire_21[13], cwire_21[14]);
fa f21_15 (pwire_21[15], swire_20[15], cwire_21[14], swire_21[14], cwire_21[15]);
fa f21_16 (pwire_21[16], swire_20[16], cwire_21[15], swire_21[15], cwire_21[16]);
fa f21_17 (pwire_21[17], swire_20[17], cwire_21[16], swire_21[16], cwire_21[17]);
fa f21_18 (pwire_21[18], swire_20[18], cwire_21[17], swire_21[17], cwire_21[18]);
fa f21_19 (pwire_21[19], swire_20[19], cwire_21[18], swire_21[18], cwire_21[19]);
fa f21_20 (pwire_21[20], swire_20[20], cwire_21[19], swire_21[19], cwire_21[20]);
fa f21_21 (pwire_21[21], swire_20[21], cwire_21[20], swire_21[20], cwire_21[21]);
fa f21_22 (pwire_21[22], swire_20[22], cwire_21[21], swire_21[21], cwire_21[22]);
fa f21_23 (pwire_21[23], swire_20[23], cwire_21[22], swire_21[22], cwire_21[23]);
fa f21_24 (pwire_21[24], swire_20[24], cwire_21[23], swire_21[23], cwire_21[24]);
fa f21_25 (pwire_21[25], swire_20[25], cwire_21[24], swire_21[24], cwire_21[25]);
fa f21_26 (pwire_21[26], swire_20[26], cwire_21[25], swire_21[25], cwire_21[26]);
fa f21_27 (pwire_21[27], swire_20[27], cwire_21[26], swire_21[26], cwire_21[27]);
fa f21_28 (pwire_21[28], swire_20[28], cwire_21[27], swire_21[27], cwire_21[28]);
fa f21_29 (pwire_21[29], swire_20[29], cwire_21[28], swire_21[28], cwire_21[29]);
fa f21_30 (pwire_21[30], swire_20[30], cwire_21[29], swire_21[29], cwire_21[30]);
fa f21_31 (pwire_21[31], swire_20[31], cwire_21[30], swire_21[30], cwire_21[31]);

//Stage21Padding
fa f21__1 (pwire_21[31], swire_20[32], cwire_21[31], swire_21[31], cwire_21[32]);
fa f21__2 (pwire_21[31], swire_20[33], cwire_21[32], swire_21[32], cwire_21[33]);
fa f21__3 (pwire_21[31], swire_20[34], cwire_21[33], swire_21[33], cwire_21[34]);
fa f21__4 (pwire_21[31], swire_20[35], cwire_21[34], swire_21[34], cwire_21[35]);
fa f21__5 (pwire_21[31], swire_20[36], cwire_21[35], swire_21[35], cwire_21[36]);
fa f21__6 (pwire_21[31], swire_20[37], cwire_21[36], swire_21[36], cwire_21[37]);
fa f21__7 (pwire_21[31], swire_20[38], cwire_21[37], swire_21[37], cwire_21[38]);
fa f21__8 (pwire_21[31], swire_20[39], cwire_21[38], swire_21[38], cwire_21[39]);
fa f21__9 (pwire_21[31], swire_20[40], cwire_21[39], swire_21[39], cwire_21[40]);
fa f21__10 (pwire_21[31], swire_20[41], cwire_21[40], swire_21[40], cwire_21[41]);
fa f21__11 (pwire_21[31], swire_20[42], cwire_21[41], swire_21[41], cwire_21[42]);

//Stage22 Partial Mul
ha f22(pwire_22[0], swire_21[0], mul[22], cwire_22[0]);
fa f22_1 (pwire_22[1], swire_21[1], cwire_22[0], swire_22[0], cwire_22[1]);
fa f22_2 (pwire_22[2], swire_21[2], cwire_22[1], swire_22[1], cwire_22[2]);
fa f22_3 (pwire_22[3], swire_21[3], cwire_22[2], swire_22[2], cwire_22[3]);
fa f22_4 (pwire_22[4], swire_21[4], cwire_22[3], swire_22[3], cwire_22[4]);
fa f22_5 (pwire_22[5], swire_21[5], cwire_22[4], swire_22[4], cwire_22[5]);
fa f22_6 (pwire_22[6], swire_21[6], cwire_22[5], swire_22[5], cwire_22[6]);
fa f22_7 (pwire_22[7], swire_21[7], cwire_22[6], swire_22[6], cwire_22[7]);
fa f22_8 (pwire_22[8], swire_21[8], cwire_22[7], swire_22[7], cwire_22[8]);
fa f22_9 (pwire_22[9], swire_21[9], cwire_22[8], swire_22[8], cwire_22[9]);
fa f22_10 (pwire_22[10], swire_21[10], cwire_22[9], swire_22[9], cwire_22[10]);
fa f22_11 (pwire_22[11], swire_21[11], cwire_22[10], swire_22[10], cwire_22[11]);
fa f22_12 (pwire_22[12], swire_21[12], cwire_22[11], swire_22[11], cwire_22[12]);
fa f22_13 (pwire_22[13], swire_21[13], cwire_22[12], swire_22[12], cwire_22[13]);
fa f22_14 (pwire_22[14], swire_21[14], cwire_22[13], swire_22[13], cwire_22[14]);
fa f22_15 (pwire_22[15], swire_21[15], cwire_22[14], swire_22[14], cwire_22[15]);
fa f22_16 (pwire_22[16], swire_21[16], cwire_22[15], swire_22[15], cwire_22[16]);
fa f22_17 (pwire_22[17], swire_21[17], cwire_22[16], swire_22[16], cwire_22[17]);
fa f22_18 (pwire_22[18], swire_21[18], cwire_22[17], swire_22[17], cwire_22[18]);
fa f22_19 (pwire_22[19], swire_21[19], cwire_22[18], swire_22[18], cwire_22[19]);
fa f22_20 (pwire_22[20], swire_21[20], cwire_22[19], swire_22[19], cwire_22[20]);
fa f22_21 (pwire_22[21], swire_21[21], cwire_22[20], swire_22[20], cwire_22[21]);
fa f22_22 (pwire_22[22], swire_21[22], cwire_22[21], swire_22[21], cwire_22[22]);
fa f22_23 (pwire_22[23], swire_21[23], cwire_22[22], swire_22[22], cwire_22[23]);
fa f22_24 (pwire_22[24], swire_21[24], cwire_22[23], swire_22[23], cwire_22[24]);
fa f22_25 (pwire_22[25], swire_21[25], cwire_22[24], swire_22[24], cwire_22[25]);
fa f22_26 (pwire_22[26], swire_21[26], cwire_22[25], swire_22[25], cwire_22[26]);
fa f22_27 (pwire_22[27], swire_21[27], cwire_22[26], swire_22[26], cwire_22[27]);
fa f22_28 (pwire_22[28], swire_21[28], cwire_22[27], swire_22[27], cwire_22[28]);
fa f22_29 (pwire_22[29], swire_21[29], cwire_22[28], swire_22[28], cwire_22[29]);
fa f22_30 (pwire_22[30], swire_21[30], cwire_22[29], swire_22[29], cwire_22[30]);
fa f22_31 (pwire_22[31], swire_21[31], cwire_22[30], swire_22[30], cwire_22[31]);

//Stage22Padding
fa f22__1 (pwire_22[31], swire_21[32], cwire_22[31], swire_22[31], cwire_22[32]);
fa f22__2 (pwire_22[31], swire_21[33], cwire_22[32], swire_22[32], cwire_22[33]);
fa f22__3 (pwire_22[31], swire_21[34], cwire_22[33], swire_22[33], cwire_22[34]);
fa f22__4 (pwire_22[31], swire_21[35], cwire_22[34], swire_22[34], cwire_22[35]);
fa f22__5 (pwire_22[31], swire_21[36], cwire_22[35], swire_22[35], cwire_22[36]);
fa f22__6 (pwire_22[31], swire_21[37], cwire_22[36], swire_22[36], cwire_22[37]);
fa f22__7 (pwire_22[31], swire_21[38], cwire_22[37], swire_22[37], cwire_22[38]);
fa f22__8 (pwire_22[31], swire_21[39], cwire_22[38], swire_22[38], cwire_22[39]);
fa f22__9 (pwire_22[31], swire_21[40], cwire_22[39], swire_22[39], cwire_22[40]);
fa f22__10 (pwire_22[31], swire_21[41], cwire_22[40], swire_22[40], cwire_22[41]);

//Stage23 Partial Mul
ha f23(pwire_23[0], swire_22[0], mul[23], cwire_23[0]);
fa f23_1 (pwire_23[1], swire_22[1], cwire_23[0], swire_23[0], cwire_23[1]);
fa f23_2 (pwire_23[2], swire_22[2], cwire_23[1], swire_23[1], cwire_23[2]);
fa f23_3 (pwire_23[3], swire_22[3], cwire_23[2], swire_23[2], cwire_23[3]);
fa f23_4 (pwire_23[4], swire_22[4], cwire_23[3], swire_23[3], cwire_23[4]);
fa f23_5 (pwire_23[5], swire_22[5], cwire_23[4], swire_23[4], cwire_23[5]);
fa f23_6 (pwire_23[6], swire_22[6], cwire_23[5], swire_23[5], cwire_23[6]);
fa f23_7 (pwire_23[7], swire_22[7], cwire_23[6], swire_23[6], cwire_23[7]);
fa f23_8 (pwire_23[8], swire_22[8], cwire_23[7], swire_23[7], cwire_23[8]);
fa f23_9 (pwire_23[9], swire_22[9], cwire_23[8], swire_23[8], cwire_23[9]);
fa f23_10 (pwire_23[10], swire_22[10], cwire_23[9], swire_23[9], cwire_23[10]);
fa f23_11 (pwire_23[11], swire_22[11], cwire_23[10], swire_23[10], cwire_23[11]);
fa f23_12 (pwire_23[12], swire_22[12], cwire_23[11], swire_23[11], cwire_23[12]);
fa f23_13 (pwire_23[13], swire_22[13], cwire_23[12], swire_23[12], cwire_23[13]);
fa f23_14 (pwire_23[14], swire_22[14], cwire_23[13], swire_23[13], cwire_23[14]);
fa f23_15 (pwire_23[15], swire_22[15], cwire_23[14], swire_23[14], cwire_23[15]);
fa f23_16 (pwire_23[16], swire_22[16], cwire_23[15], swire_23[15], cwire_23[16]);
fa f23_17 (pwire_23[17], swire_22[17], cwire_23[16], swire_23[16], cwire_23[17]);
fa f23_18 (pwire_23[18], swire_22[18], cwire_23[17], swire_23[17], cwire_23[18]);
fa f23_19 (pwire_23[19], swire_22[19], cwire_23[18], swire_23[18], cwire_23[19]);
fa f23_20 (pwire_23[20], swire_22[20], cwire_23[19], swire_23[19], cwire_23[20]);
fa f23_21 (pwire_23[21], swire_22[21], cwire_23[20], swire_23[20], cwire_23[21]);
fa f23_22 (pwire_23[22], swire_22[22], cwire_23[21], swire_23[21], cwire_23[22]);
fa f23_23 (pwire_23[23], swire_22[23], cwire_23[22], swire_23[22], cwire_23[23]);
fa f23_24 (pwire_23[24], swire_22[24], cwire_23[23], swire_23[23], cwire_23[24]);
fa f23_25 (pwire_23[25], swire_22[25], cwire_23[24], swire_23[24], cwire_23[25]);
fa f23_26 (pwire_23[26], swire_22[26], cwire_23[25], swire_23[25], cwire_23[26]);
fa f23_27 (pwire_23[27], swire_22[27], cwire_23[26], swire_23[26], cwire_23[27]);
fa f23_28 (pwire_23[28], swire_22[28], cwire_23[27], swire_23[27], cwire_23[28]);
fa f23_29 (pwire_23[29], swire_22[29], cwire_23[28], swire_23[28], cwire_23[29]);
fa f23_30 (pwire_23[30], swire_22[30], cwire_23[29], swire_23[29], cwire_23[30]);
fa f23_31 (pwire_23[31], swire_22[31], cwire_23[30], swire_23[30], cwire_23[31]);

//Stage23Padding
fa f23__1 (pwire_23[31], swire_22[32], cwire_23[31], swire_23[31], cwire_23[32]);
fa f23__2 (pwire_23[31], swire_22[33], cwire_23[32], swire_23[32], cwire_23[33]);
fa f23__3 (pwire_23[31], swire_22[34], cwire_23[33], swire_23[33], cwire_23[34]);
fa f23__4 (pwire_23[31], swire_22[35], cwire_23[34], swire_23[34], cwire_23[35]);
fa f23__5 (pwire_23[31], swire_22[36], cwire_23[35], swire_23[35], cwire_23[36]);
fa f23__6 (pwire_23[31], swire_22[37], cwire_23[36], swire_23[36], cwire_23[37]);
fa f23__7 (pwire_23[31], swire_22[38], cwire_23[37], swire_23[37], cwire_23[38]);
fa f23__8 (pwire_23[31], swire_22[39], cwire_23[38], swire_23[38], cwire_23[39]);
fa f23__9 (pwire_23[31], swire_22[40], cwire_23[39], swire_23[39], cwire_23[40]);

//Stage24 Partial Mul
ha f24(pwire_24[0], swire_23[0], mul[24], cwire_24[0]);
fa f24_1 (pwire_24[1], swire_23[1], cwire_24[0], swire_24[0], cwire_24[1]);
fa f24_2 (pwire_24[2], swire_23[2], cwire_24[1], swire_24[1], cwire_24[2]);
fa f24_3 (pwire_24[3], swire_23[3], cwire_24[2], swire_24[2], cwire_24[3]);
fa f24_4 (pwire_24[4], swire_23[4], cwire_24[3], swire_24[3], cwire_24[4]);
fa f24_5 (pwire_24[5], swire_23[5], cwire_24[4], swire_24[4], cwire_24[5]);
fa f24_6 (pwire_24[6], swire_23[6], cwire_24[5], swire_24[5], cwire_24[6]);
fa f24_7 (pwire_24[7], swire_23[7], cwire_24[6], swire_24[6], cwire_24[7]);
fa f24_8 (pwire_24[8], swire_23[8], cwire_24[7], swire_24[7], cwire_24[8]);
fa f24_9 (pwire_24[9], swire_23[9], cwire_24[8], swire_24[8], cwire_24[9]);
fa f24_10 (pwire_24[10], swire_23[10], cwire_24[9], swire_24[9], cwire_24[10]);
fa f24_11 (pwire_24[11], swire_23[11], cwire_24[10], swire_24[10], cwire_24[11]);
fa f24_12 (pwire_24[12], swire_23[12], cwire_24[11], swire_24[11], cwire_24[12]);
fa f24_13 (pwire_24[13], swire_23[13], cwire_24[12], swire_24[12], cwire_24[13]);
fa f24_14 (pwire_24[14], swire_23[14], cwire_24[13], swire_24[13], cwire_24[14]);
fa f24_15 (pwire_24[15], swire_23[15], cwire_24[14], swire_24[14], cwire_24[15]);
fa f24_16 (pwire_24[16], swire_23[16], cwire_24[15], swire_24[15], cwire_24[16]);
fa f24_17 (pwire_24[17], swire_23[17], cwire_24[16], swire_24[16], cwire_24[17]);
fa f24_18 (pwire_24[18], swire_23[18], cwire_24[17], swire_24[17], cwire_24[18]);
fa f24_19 (pwire_24[19], swire_23[19], cwire_24[18], swire_24[18], cwire_24[19]);
fa f24_20 (pwire_24[20], swire_23[20], cwire_24[19], swire_24[19], cwire_24[20]);
fa f24_21 (pwire_24[21], swire_23[21], cwire_24[20], swire_24[20], cwire_24[21]);
fa f24_22 (pwire_24[22], swire_23[22], cwire_24[21], swire_24[21], cwire_24[22]);
fa f24_23 (pwire_24[23], swire_23[23], cwire_24[22], swire_24[22], cwire_24[23]);
fa f24_24 (pwire_24[24], swire_23[24], cwire_24[23], swire_24[23], cwire_24[24]);
fa f24_25 (pwire_24[25], swire_23[25], cwire_24[24], swire_24[24], cwire_24[25]);
fa f24_26 (pwire_24[26], swire_23[26], cwire_24[25], swire_24[25], cwire_24[26]);
fa f24_27 (pwire_24[27], swire_23[27], cwire_24[26], swire_24[26], cwire_24[27]);
fa f24_28 (pwire_24[28], swire_23[28], cwire_24[27], swire_24[27], cwire_24[28]);
fa f24_29 (pwire_24[29], swire_23[29], cwire_24[28], swire_24[28], cwire_24[29]);
fa f24_30 (pwire_24[30], swire_23[30], cwire_24[29], swire_24[29], cwire_24[30]);
fa f24_31 (pwire_24[31], swire_23[31], cwire_24[30], swire_24[30], cwire_24[31]);

//Stage24Padding
fa f24__1 (pwire_24[31], swire_23[32], cwire_24[31], swire_24[31], cwire_24[32]);
fa f24__2 (pwire_24[31], swire_23[33], cwire_24[32], swire_24[32], cwire_24[33]);
fa f24__3 (pwire_24[31], swire_23[34], cwire_24[33], swire_24[33], cwire_24[34]);
fa f24__4 (pwire_24[31], swire_23[35], cwire_24[34], swire_24[34], cwire_24[35]);
fa f24__5 (pwire_24[31], swire_23[36], cwire_24[35], swire_24[35], cwire_24[36]);
fa f24__6 (pwire_24[31], swire_23[37], cwire_24[36], swire_24[36], cwire_24[37]);
fa f24__7 (pwire_24[31], swire_23[38], cwire_24[37], swire_24[37], cwire_24[38]);
fa f24__8 (pwire_24[31], swire_23[39], cwire_24[38], swire_24[38], cwire_24[39]);

//Stage25 Partial Mul
ha f25(pwire_25[0], swire_24[0], mul[25], cwire_25[0]);
fa f25_1 (pwire_25[1], swire_24[1], cwire_25[0], swire_25[0], cwire_25[1]);
fa f25_2 (pwire_25[2], swire_24[2], cwire_25[1], swire_25[1], cwire_25[2]);
fa f25_3 (pwire_25[3], swire_24[3], cwire_25[2], swire_25[2], cwire_25[3]);
fa f25_4 (pwire_25[4], swire_24[4], cwire_25[3], swire_25[3], cwire_25[4]);
fa f25_5 (pwire_25[5], swire_24[5], cwire_25[4], swire_25[4], cwire_25[5]);
fa f25_6 (pwire_25[6], swire_24[6], cwire_25[5], swire_25[5], cwire_25[6]);
fa f25_7 (pwire_25[7], swire_24[7], cwire_25[6], swire_25[6], cwire_25[7]);
fa f25_8 (pwire_25[8], swire_24[8], cwire_25[7], swire_25[7], cwire_25[8]);
fa f25_9 (pwire_25[9], swire_24[9], cwire_25[8], swire_25[8], cwire_25[9]);
fa f25_10 (pwire_25[10], swire_24[10], cwire_25[9], swire_25[9], cwire_25[10]);
fa f25_11 (pwire_25[11], swire_24[11], cwire_25[10], swire_25[10], cwire_25[11]);
fa f25_12 (pwire_25[12], swire_24[12], cwire_25[11], swire_25[11], cwire_25[12]);
fa f25_13 (pwire_25[13], swire_24[13], cwire_25[12], swire_25[12], cwire_25[13]);
fa f25_14 (pwire_25[14], swire_24[14], cwire_25[13], swire_25[13], cwire_25[14]);
fa f25_15 (pwire_25[15], swire_24[15], cwire_25[14], swire_25[14], cwire_25[15]);
fa f25_16 (pwire_25[16], swire_24[16], cwire_25[15], swire_25[15], cwire_25[16]);
fa f25_17 (pwire_25[17], swire_24[17], cwire_25[16], swire_25[16], cwire_25[17]);
fa f25_18 (pwire_25[18], swire_24[18], cwire_25[17], swire_25[17], cwire_25[18]);
fa f25_19 (pwire_25[19], swire_24[19], cwire_25[18], swire_25[18], cwire_25[19]);
fa f25_20 (pwire_25[20], swire_24[20], cwire_25[19], swire_25[19], cwire_25[20]);
fa f25_21 (pwire_25[21], swire_24[21], cwire_25[20], swire_25[20], cwire_25[21]);
fa f25_22 (pwire_25[22], swire_24[22], cwire_25[21], swire_25[21], cwire_25[22]);
fa f25_23 (pwire_25[23], swire_24[23], cwire_25[22], swire_25[22], cwire_25[23]);
fa f25_24 (pwire_25[24], swire_24[24], cwire_25[23], swire_25[23], cwire_25[24]);
fa f25_25 (pwire_25[25], swire_24[25], cwire_25[24], swire_25[24], cwire_25[25]);
fa f25_26 (pwire_25[26], swire_24[26], cwire_25[25], swire_25[25], cwire_25[26]);
fa f25_27 (pwire_25[27], swire_24[27], cwire_25[26], swire_25[26], cwire_25[27]);
fa f25_28 (pwire_25[28], swire_24[28], cwire_25[27], swire_25[27], cwire_25[28]);
fa f25_29 (pwire_25[29], swire_24[29], cwire_25[28], swire_25[28], cwire_25[29]);
fa f25_30 (pwire_25[30], swire_24[30], cwire_25[29], swire_25[29], cwire_25[30]);
fa f25_31 (pwire_25[31], swire_24[31], cwire_25[30], swire_25[30], cwire_25[31]);

//Stage25Padding
fa f25__1 (pwire_25[31], swire_24[32], cwire_25[31], swire_25[31], cwire_25[32]);
fa f25__2 (pwire_25[31], swire_24[33], cwire_25[32], swire_25[32], cwire_25[33]);
fa f25__3 (pwire_25[31], swire_24[34], cwire_25[33], swire_25[33], cwire_25[34]);
fa f25__4 (pwire_25[31], swire_24[35], cwire_25[34], swire_25[34], cwire_25[35]);
fa f25__5 (pwire_25[31], swire_24[36], cwire_25[35], swire_25[35], cwire_25[36]);
fa f25__6 (pwire_25[31], swire_24[37], cwire_25[36], swire_25[36], cwire_25[37]);
fa f25__7 (pwire_25[31], swire_24[38], cwire_25[37], swire_25[37], cwire_25[38]);

//Stage26 Partial Mul
ha f26(pwire_26[0], swire_25[0], mul[26], cwire_26[0]);
fa f26_1 (pwire_26[1], swire_25[1], cwire_26[0], swire_26[0], cwire_26[1]);
fa f26_2 (pwire_26[2], swire_25[2], cwire_26[1], swire_26[1], cwire_26[2]);
fa f26_3 (pwire_26[3], swire_25[3], cwire_26[2], swire_26[2], cwire_26[3]);
fa f26_4 (pwire_26[4], swire_25[4], cwire_26[3], swire_26[3], cwire_26[4]);
fa f26_5 (pwire_26[5], swire_25[5], cwire_26[4], swire_26[4], cwire_26[5]);
fa f26_6 (pwire_26[6], swire_25[6], cwire_26[5], swire_26[5], cwire_26[6]);
fa f26_7 (pwire_26[7], swire_25[7], cwire_26[6], swire_26[6], cwire_26[7]);
fa f26_8 (pwire_26[8], swire_25[8], cwire_26[7], swire_26[7], cwire_26[8]);
fa f26_9 (pwire_26[9], swire_25[9], cwire_26[8], swire_26[8], cwire_26[9]);
fa f26_10 (pwire_26[10], swire_25[10], cwire_26[9], swire_26[9], cwire_26[10]);
fa f26_11 (pwire_26[11], swire_25[11], cwire_26[10], swire_26[10], cwire_26[11]);
fa f26_12 (pwire_26[12], swire_25[12], cwire_26[11], swire_26[11], cwire_26[12]);
fa f26_13 (pwire_26[13], swire_25[13], cwire_26[12], swire_26[12], cwire_26[13]);
fa f26_14 (pwire_26[14], swire_25[14], cwire_26[13], swire_26[13], cwire_26[14]);
fa f26_15 (pwire_26[15], swire_25[15], cwire_26[14], swire_26[14], cwire_26[15]);
fa f26_16 (pwire_26[16], swire_25[16], cwire_26[15], swire_26[15], cwire_26[16]);
fa f26_17 (pwire_26[17], swire_25[17], cwire_26[16], swire_26[16], cwire_26[17]);
fa f26_18 (pwire_26[18], swire_25[18], cwire_26[17], swire_26[17], cwire_26[18]);
fa f26_19 (pwire_26[19], swire_25[19], cwire_26[18], swire_26[18], cwire_26[19]);
fa f26_20 (pwire_26[20], swire_25[20], cwire_26[19], swire_26[19], cwire_26[20]);
fa f26_21 (pwire_26[21], swire_25[21], cwire_26[20], swire_26[20], cwire_26[21]);
fa f26_22 (pwire_26[22], swire_25[22], cwire_26[21], swire_26[21], cwire_26[22]);
fa f26_23 (pwire_26[23], swire_25[23], cwire_26[22], swire_26[22], cwire_26[23]);
fa f26_24 (pwire_26[24], swire_25[24], cwire_26[23], swire_26[23], cwire_26[24]);
fa f26_25 (pwire_26[25], swire_25[25], cwire_26[24], swire_26[24], cwire_26[25]);
fa f26_26 (pwire_26[26], swire_25[26], cwire_26[25], swire_26[25], cwire_26[26]);
fa f26_27 (pwire_26[27], swire_25[27], cwire_26[26], swire_26[26], cwire_26[27]);
fa f26_28 (pwire_26[28], swire_25[28], cwire_26[27], swire_26[27], cwire_26[28]);
fa f26_29 (pwire_26[29], swire_25[29], cwire_26[28], swire_26[28], cwire_26[29]);
fa f26_30 (pwire_26[30], swire_25[30], cwire_26[29], swire_26[29], cwire_26[30]);
fa f26_31 (pwire_26[31], swire_25[31], cwire_26[30], swire_26[30], cwire_26[31]);

//Stage26Padding
fa f26__1 (pwire_26[31], swire_25[32], cwire_26[31], swire_26[31], cwire_26[32]);
fa f26__2 (pwire_26[31], swire_25[33], cwire_26[32], swire_26[32], cwire_26[33]);
fa f26__3 (pwire_26[31], swire_25[34], cwire_26[33], swire_26[33], cwire_26[34]);
fa f26__4 (pwire_26[31], swire_25[35], cwire_26[34], swire_26[34], cwire_26[35]);
fa f26__5 (pwire_26[31], swire_25[36], cwire_26[35], swire_26[35], cwire_26[36]);
fa f26__6 (pwire_26[31], swire_25[37], cwire_26[36], swire_26[36], cwire_26[37]);

//Stage27 Partial Mul
ha f27(pwire_27[0], swire_26[0], mul[27], cwire_27[0]);
fa f27_1 (pwire_27[1], swire_26[1], cwire_27[0], swire_27[0], cwire_27[1]);
fa f27_2 (pwire_27[2], swire_26[2], cwire_27[1], swire_27[1], cwire_27[2]);
fa f27_3 (pwire_27[3], swire_26[3], cwire_27[2], swire_27[2], cwire_27[3]);
fa f27_4 (pwire_27[4], swire_26[4], cwire_27[3], swire_27[3], cwire_27[4]);
fa f27_5 (pwire_27[5], swire_26[5], cwire_27[4], swire_27[4], cwire_27[5]);
fa f27_6 (pwire_27[6], swire_26[6], cwire_27[5], swire_27[5], cwire_27[6]);
fa f27_7 (pwire_27[7], swire_26[7], cwire_27[6], swire_27[6], cwire_27[7]);
fa f27_8 (pwire_27[8], swire_26[8], cwire_27[7], swire_27[7], cwire_27[8]);
fa f27_9 (pwire_27[9], swire_26[9], cwire_27[8], swire_27[8], cwire_27[9]);
fa f27_10 (pwire_27[10], swire_26[10], cwire_27[9], swire_27[9], cwire_27[10]);
fa f27_11 (pwire_27[11], swire_26[11], cwire_27[10], swire_27[10], cwire_27[11]);
fa f27_12 (pwire_27[12], swire_26[12], cwire_27[11], swire_27[11], cwire_27[12]);
fa f27_13 (pwire_27[13], swire_26[13], cwire_27[12], swire_27[12], cwire_27[13]);
fa f27_14 (pwire_27[14], swire_26[14], cwire_27[13], swire_27[13], cwire_27[14]);
fa f27_15 (pwire_27[15], swire_26[15], cwire_27[14], swire_27[14], cwire_27[15]);
fa f27_16 (pwire_27[16], swire_26[16], cwire_27[15], swire_27[15], cwire_27[16]);
fa f27_17 (pwire_27[17], swire_26[17], cwire_27[16], swire_27[16], cwire_27[17]);
fa f27_18 (pwire_27[18], swire_26[18], cwire_27[17], swire_27[17], cwire_27[18]);
fa f27_19 (pwire_27[19], swire_26[19], cwire_27[18], swire_27[18], cwire_27[19]);
fa f27_20 (pwire_27[20], swire_26[20], cwire_27[19], swire_27[19], cwire_27[20]);
fa f27_21 (pwire_27[21], swire_26[21], cwire_27[20], swire_27[20], cwire_27[21]);
fa f27_22 (pwire_27[22], swire_26[22], cwire_27[21], swire_27[21], cwire_27[22]);
fa f27_23 (pwire_27[23], swire_26[23], cwire_27[22], swire_27[22], cwire_27[23]);
fa f27_24 (pwire_27[24], swire_26[24], cwire_27[23], swire_27[23], cwire_27[24]);
fa f27_25 (pwire_27[25], swire_26[25], cwire_27[24], swire_27[24], cwire_27[25]);
fa f27_26 (pwire_27[26], swire_26[26], cwire_27[25], swire_27[25], cwire_27[26]);
fa f27_27 (pwire_27[27], swire_26[27], cwire_27[26], swire_27[26], cwire_27[27]);
fa f27_28 (pwire_27[28], swire_26[28], cwire_27[27], swire_27[27], cwire_27[28]);
fa f27_29 (pwire_27[29], swire_26[29], cwire_27[28], swire_27[28], cwire_27[29]);
fa f27_30 (pwire_27[30], swire_26[30], cwire_27[29], swire_27[29], cwire_27[30]);
fa f27_31 (pwire_27[31], swire_26[31], cwire_27[30], swire_27[30], cwire_27[31]);

//Stage27Padding
fa f27__1 (pwire_27[31], swire_26[32], cwire_27[31], swire_27[31], cwire_27[32]);
fa f27__2 (pwire_27[31], swire_26[33], cwire_27[32], swire_27[32], cwire_27[33]);
fa f27__3 (pwire_27[31], swire_26[34], cwire_27[33], swire_27[33], cwire_27[34]);
fa f27__4 (pwire_27[31], swire_26[35], cwire_27[34], swire_27[34], cwire_27[35]);
fa f27__5 (pwire_27[31], swire_26[36], cwire_27[35], swire_27[35], cwire_27[36]);

//Stage28 Partial Mul
ha f28(pwire_28[0], swire_27[0], mul[28], cwire_28[0]);
fa f28_1 (pwire_28[1], swire_27[1], cwire_28[0], swire_28[0], cwire_28[1]);
fa f28_2 (pwire_28[2], swire_27[2], cwire_28[1], swire_28[1], cwire_28[2]);
fa f28_3 (pwire_28[3], swire_27[3], cwire_28[2], swire_28[2], cwire_28[3]);
fa f28_4 (pwire_28[4], swire_27[4], cwire_28[3], swire_28[3], cwire_28[4]);
fa f28_5 (pwire_28[5], swire_27[5], cwire_28[4], swire_28[4], cwire_28[5]);
fa f28_6 (pwire_28[6], swire_27[6], cwire_28[5], swire_28[5], cwire_28[6]);
fa f28_7 (pwire_28[7], swire_27[7], cwire_28[6], swire_28[6], cwire_28[7]);
fa f28_8 (pwire_28[8], swire_27[8], cwire_28[7], swire_28[7], cwire_28[8]);
fa f28_9 (pwire_28[9], swire_27[9], cwire_28[8], swire_28[8], cwire_28[9]);
fa f28_10 (pwire_28[10], swire_27[10], cwire_28[9], swire_28[9], cwire_28[10]);
fa f28_11 (pwire_28[11], swire_27[11], cwire_28[10], swire_28[10], cwire_28[11]);
fa f28_12 (pwire_28[12], swire_27[12], cwire_28[11], swire_28[11], cwire_28[12]);
fa f28_13 (pwire_28[13], swire_27[13], cwire_28[12], swire_28[12], cwire_28[13]);
fa f28_14 (pwire_28[14], swire_27[14], cwire_28[13], swire_28[13], cwire_28[14]);
fa f28_15 (pwire_28[15], swire_27[15], cwire_28[14], swire_28[14], cwire_28[15]);
fa f28_16 (pwire_28[16], swire_27[16], cwire_28[15], swire_28[15], cwire_28[16]);
fa f28_17 (pwire_28[17], swire_27[17], cwire_28[16], swire_28[16], cwire_28[17]);
fa f28_18 (pwire_28[18], swire_27[18], cwire_28[17], swire_28[17], cwire_28[18]);
fa f28_19 (pwire_28[19], swire_27[19], cwire_28[18], swire_28[18], cwire_28[19]);
fa f28_20 (pwire_28[20], swire_27[20], cwire_28[19], swire_28[19], cwire_28[20]);
fa f28_21 (pwire_28[21], swire_27[21], cwire_28[20], swire_28[20], cwire_28[21]);
fa f28_22 (pwire_28[22], swire_27[22], cwire_28[21], swire_28[21], cwire_28[22]);
fa f28_23 (pwire_28[23], swire_27[23], cwire_28[22], swire_28[22], cwire_28[23]);
fa f28_24 (pwire_28[24], swire_27[24], cwire_28[23], swire_28[23], cwire_28[24]);
fa f28_25 (pwire_28[25], swire_27[25], cwire_28[24], swire_28[24], cwire_28[25]);
fa f28_26 (pwire_28[26], swire_27[26], cwire_28[25], swire_28[25], cwire_28[26]);
fa f28_27 (pwire_28[27], swire_27[27], cwire_28[26], swire_28[26], cwire_28[27]);
fa f28_28 (pwire_28[28], swire_27[28], cwire_28[27], swire_28[27], cwire_28[28]);
fa f28_29 (pwire_28[29], swire_27[29], cwire_28[28], swire_28[28], cwire_28[29]);
fa f28_30 (pwire_28[30], swire_27[30], cwire_28[29], swire_28[29], cwire_28[30]);
fa f28_31 (pwire_28[31], swire_27[31], cwire_28[30], swire_28[30], cwire_28[31]);

//Stage28Padding
fa f28__1 (pwire_28[31], swire_27[32], cwire_28[31], swire_28[31], cwire_28[32]);
fa f28__2 (pwire_28[31], swire_27[33], cwire_28[32], swire_28[32], cwire_28[33]);
fa f28__3 (pwire_28[31], swire_27[34], cwire_28[33], swire_28[33], cwire_28[34]);
fa f28__4 (pwire_28[31], swire_27[35], cwire_28[34], swire_28[34], cwire_28[35]);

//Stage29 Partial Mul
ha f29(pwire_29[0], swire_28[0], mul[29], cwire_29[0]);
fa f29_1 (pwire_29[1], swire_28[1], cwire_29[0], swire_29[0], cwire_29[1]);
fa f29_2 (pwire_29[2], swire_28[2], cwire_29[1], swire_29[1], cwire_29[2]);
fa f29_3 (pwire_29[3], swire_28[3], cwire_29[2], swire_29[2], cwire_29[3]);
fa f29_4 (pwire_29[4], swire_28[4], cwire_29[3], swire_29[3], cwire_29[4]);
fa f29_5 (pwire_29[5], swire_28[5], cwire_29[4], swire_29[4], cwire_29[5]);
fa f29_6 (pwire_29[6], swire_28[6], cwire_29[5], swire_29[5], cwire_29[6]);
fa f29_7 (pwire_29[7], swire_28[7], cwire_29[6], swire_29[6], cwire_29[7]);
fa f29_8 (pwire_29[8], swire_28[8], cwire_29[7], swire_29[7], cwire_29[8]);
fa f29_9 (pwire_29[9], swire_28[9], cwire_29[8], swire_29[8], cwire_29[9]);
fa f29_10 (pwire_29[10], swire_28[10], cwire_29[9], swire_29[9], cwire_29[10]);
fa f29_11 (pwire_29[11], swire_28[11], cwire_29[10], swire_29[10], cwire_29[11]);
fa f29_12 (pwire_29[12], swire_28[12], cwire_29[11], swire_29[11], cwire_29[12]);
fa f29_13 (pwire_29[13], swire_28[13], cwire_29[12], swire_29[12], cwire_29[13]);
fa f29_14 (pwire_29[14], swire_28[14], cwire_29[13], swire_29[13], cwire_29[14]);
fa f29_15 (pwire_29[15], swire_28[15], cwire_29[14], swire_29[14], cwire_29[15]);
fa f29_16 (pwire_29[16], swire_28[16], cwire_29[15], swire_29[15], cwire_29[16]);
fa f29_17 (pwire_29[17], swire_28[17], cwire_29[16], swire_29[16], cwire_29[17]);
fa f29_18 (pwire_29[18], swire_28[18], cwire_29[17], swire_29[17], cwire_29[18]);
fa f29_19 (pwire_29[19], swire_28[19], cwire_29[18], swire_29[18], cwire_29[19]);
fa f29_20 (pwire_29[20], swire_28[20], cwire_29[19], swire_29[19], cwire_29[20]);
fa f29_21 (pwire_29[21], swire_28[21], cwire_29[20], swire_29[20], cwire_29[21]);
fa f29_22 (pwire_29[22], swire_28[22], cwire_29[21], swire_29[21], cwire_29[22]);
fa f29_23 (pwire_29[23], swire_28[23], cwire_29[22], swire_29[22], cwire_29[23]);
fa f29_24 (pwire_29[24], swire_28[24], cwire_29[23], swire_29[23], cwire_29[24]);
fa f29_25 (pwire_29[25], swire_28[25], cwire_29[24], swire_29[24], cwire_29[25]);
fa f29_26 (pwire_29[26], swire_28[26], cwire_29[25], swire_29[25], cwire_29[26]);
fa f29_27 (pwire_29[27], swire_28[27], cwire_29[26], swire_29[26], cwire_29[27]);
fa f29_28 (pwire_29[28], swire_28[28], cwire_29[27], swire_29[27], cwire_29[28]);
fa f29_29 (pwire_29[29], swire_28[29], cwire_29[28], swire_29[28], cwire_29[29]);
fa f29_30 (pwire_29[30], swire_28[30], cwire_29[29], swire_29[29], cwire_29[30]);
fa f29_31 (pwire_29[31], swire_28[31], cwire_29[30], swire_29[30], cwire_29[31]);

//Stage29Padding
fa f29__1 (pwire_29[31], swire_28[32], cwire_29[31], swire_29[31], cwire_29[32]);
fa f29__2 (pwire_29[31], swire_28[33], cwire_29[32], swire_29[32], cwire_29[33]);
fa f29__3 (pwire_29[31], swire_28[34], cwire_29[33], swire_29[33], cwire_29[34]);

//Stage30 Partial Mul
ha f30(pwire_30[0], swire_29[0], mul[30], cwire_30[0]);
fa f30_1 (pwire_30[1], swire_29[1], cwire_30[0], swire_30[0], cwire_30[1]);
fa f30_2 (pwire_30[2], swire_29[2], cwire_30[1], swire_30[1], cwire_30[2]);
fa f30_3 (pwire_30[3], swire_29[3], cwire_30[2], swire_30[2], cwire_30[3]);
fa f30_4 (pwire_30[4], swire_29[4], cwire_30[3], swire_30[3], cwire_30[4]);
fa f30_5 (pwire_30[5], swire_29[5], cwire_30[4], swire_30[4], cwire_30[5]);
fa f30_6 (pwire_30[6], swire_29[6], cwire_30[5], swire_30[5], cwire_30[6]);
fa f30_7 (pwire_30[7], swire_29[7], cwire_30[6], swire_30[6], cwire_30[7]);
fa f30_8 (pwire_30[8], swire_29[8], cwire_30[7], swire_30[7], cwire_30[8]);
fa f30_9 (pwire_30[9], swire_29[9], cwire_30[8], swire_30[8], cwire_30[9]);
fa f30_10 (pwire_30[10], swire_29[10], cwire_30[9], swire_30[9], cwire_30[10]);
fa f30_11 (pwire_30[11], swire_29[11], cwire_30[10], swire_30[10], cwire_30[11]);
fa f30_12 (pwire_30[12], swire_29[12], cwire_30[11], swire_30[11], cwire_30[12]);
fa f30_13 (pwire_30[13], swire_29[13], cwire_30[12], swire_30[12], cwire_30[13]);
fa f30_14 (pwire_30[14], swire_29[14], cwire_30[13], swire_30[13], cwire_30[14]);
fa f30_15 (pwire_30[15], swire_29[15], cwire_30[14], swire_30[14], cwire_30[15]);
fa f30_16 (pwire_30[16], swire_29[16], cwire_30[15], swire_30[15], cwire_30[16]);
fa f30_17 (pwire_30[17], swire_29[17], cwire_30[16], swire_30[16], cwire_30[17]);
fa f30_18 (pwire_30[18], swire_29[18], cwire_30[17], swire_30[17], cwire_30[18]);
fa f30_19 (pwire_30[19], swire_29[19], cwire_30[18], swire_30[18], cwire_30[19]);
fa f30_20 (pwire_30[20], swire_29[20], cwire_30[19], swire_30[19], cwire_30[20]);
fa f30_21 (pwire_30[21], swire_29[21], cwire_30[20], swire_30[20], cwire_30[21]);
fa f30_22 (pwire_30[22], swire_29[22], cwire_30[21], swire_30[21], cwire_30[22]);
fa f30_23 (pwire_30[23], swire_29[23], cwire_30[22], swire_30[22], cwire_30[23]);
fa f30_24 (pwire_30[24], swire_29[24], cwire_30[23], swire_30[23], cwire_30[24]);
fa f30_25 (pwire_30[25], swire_29[25], cwire_30[24], swire_30[24], cwire_30[25]);
fa f30_26 (pwire_30[26], swire_29[26], cwire_30[25], swire_30[25], cwire_30[26]);
fa f30_27 (pwire_30[27], swire_29[27], cwire_30[26], swire_30[26], cwire_30[27]);
fa f30_28 (pwire_30[28], swire_29[28], cwire_30[27], swire_30[27], cwire_30[28]);
fa f30_29 (pwire_30[29], swire_29[29], cwire_30[28], swire_30[28], cwire_30[29]);
fa f30_30 (pwire_30[30], swire_29[30], cwire_30[29], swire_30[29], cwire_30[30]);
fa f30_31 (pwire_30[31], swire_29[31], cwire_30[30], swire_30[30], cwire_30[31]);

//Stage30Padding
fa f30__1 (pwire_30[31], swire_29[32], cwire_30[31], swire_30[31], cwire_30[32]);
fa f30__2 (pwire_30[31], swire_29[33], cwire_30[32], swire_30[32], cwire_30[33]);

//Stage31 Partial Mul
fa f31(pwire_31[0], swire_30[0], b[31], mul[31], cwire_31[0]);
fa f31_1 (pwire_31[1], swire_30[1], cwire_31[0], mul[32], cwire_31[1]);
fa f31_2 (pwire_31[2], swire_30[2], cwire_31[1], mul[33], cwire_31[2]);
fa f31_3 (pwire_31[3], swire_30[3], cwire_31[2], mul[34], cwire_31[3]);
fa f31_4 (pwire_31[4], swire_30[4], cwire_31[3], mul[35], cwire_31[4]);
fa f31_5 (pwire_31[5], swire_30[5], cwire_31[4], mul[36], cwire_31[5]);
fa f31_6 (pwire_31[6], swire_30[6], cwire_31[5], mul[37], cwire_31[6]);
fa f31_7 (pwire_31[7], swire_30[7], cwire_31[6], mul[38], cwire_31[7]);
fa f31_8 (pwire_31[8], swire_30[8], cwire_31[7], mul[39], cwire_31[8]);
fa f31_9 (pwire_31[9], swire_30[9], cwire_31[8], mul[40], cwire_31[9]);
fa f31_10 (pwire_31[10], swire_30[10], cwire_31[9], mul[41], cwire_31[10]);
fa f31_11 (pwire_31[11], swire_30[11], cwire_31[10], mul[42], cwire_31[11]);
fa f31_12 (pwire_31[12], swire_30[12], cwire_31[11], mul[43], cwire_31[12]);
fa f31_13 (pwire_31[13], swire_30[13], cwire_31[12], mul[44], cwire_31[13]);
fa f31_14 (pwire_31[14], swire_30[14], cwire_31[13], mul[45], cwire_31[14]);
fa f31_15 (pwire_31[15], swire_30[15], cwire_31[14], mul[46], cwire_31[15]);
fa f31_16 (pwire_31[16], swire_30[16], cwire_31[15], mul[47], cwire_31[16]);
fa f31_17 (pwire_31[17], swire_30[17], cwire_31[16], mul[48], cwire_31[17]);
fa f31_18 (pwire_31[18], swire_30[18], cwire_31[17], mul[49], cwire_31[18]);
fa f31_19 (pwire_31[19], swire_30[19], cwire_31[18], mul[50], cwire_31[19]);
fa f31_20 (pwire_31[20], swire_30[20], cwire_31[19], mul[51], cwire_31[20]);
fa f31_21 (pwire_31[21], swire_30[21], cwire_31[20], mul[52], cwire_31[21]);
fa f31_22 (pwire_31[22], swire_30[22], cwire_31[21], mul[53], cwire_31[22]);
fa f31_23 (pwire_31[23], swire_30[23], cwire_31[22], mul[54], cwire_31[23]);
fa f31_24 (pwire_31[24], swire_30[24], cwire_31[23], mul[55], cwire_31[24]);
fa f31_25 (pwire_31[25], swire_30[25], cwire_31[24], mul[56], cwire_31[25]);
fa f31_26 (pwire_31[26], swire_30[26], cwire_31[25], mul[57], cwire_31[26]);
fa f31_27 (pwire_31[27], swire_30[27], cwire_31[26], mul[58], cwire_31[27]);
fa f31_28 (pwire_31[28], swire_30[28], cwire_31[27], mul[59], cwire_31[28]);
fa f31_29 (pwire_31[29], swire_30[29], cwire_31[28], mul[60], cwire_31[29]);
fa f31_30 (pwire_31[30], swire_30[30], cwire_31[29], mul[61], cwire_31[30]);
fa f31_31 (pwire_31[31], swire_30[31], cwire_31[30], mul[62], cwire_31[31]);

//Stage31Padding
fa f31__1 (pwire_31[31], swire_30[32], cwire_31[31], mul[63], cwire_31[32]);

assign mul[0] = a[0] & b[0];
assign pwire_0 = b[0] ? a : 0;
assign pwire_1 = b[1] ? a : 0;
assign pwire_2 = b[2] ? a : 0;
assign pwire_3 = b[3] ? a : 0;
assign pwire_4 = b[4] ? a : 0;
assign pwire_5 = b[5] ? a : 0;
assign pwire_6 = b[6] ? a : 0;
assign pwire_7 = b[7] ? a : 0;
assign pwire_8 = b[8] ? a : 0;
assign pwire_9 = b[9] ? a : 0;
assign pwire_10 = b[10] ? a : 0;
assign pwire_11 = b[11] ? a : 0;
assign pwire_12 = b[12] ? a : 0;
assign pwire_13 = b[13] ? a : 0;
assign pwire_14 = b[14] ? a : 0;
assign pwire_15 = b[15] ? a : 0;
assign pwire_16 = b[16] ? a : 0;
assign pwire_17 = b[17] ? a : 0;
assign pwire_18 = b[18] ? a : 0;
assign pwire_19 = b[19] ? a : 0;
assign pwire_20 = b[20] ? a : 0;
assign pwire_21 = b[21] ? a : 0;
assign pwire_22 = b[22] ? a : 0;
assign pwire_23 = b[23] ? a : 0;
assign pwire_24 = b[24] ? a : 0;
assign pwire_25 = b[25] ? a : 0;
assign pwire_26 = b[26] ? a : 0;
assign pwire_27 = b[27] ? a : 0;
assign pwire_28 = b[28] ? a : 0;
assign pwire_29 = b[29] ? a : 0;
assign pwire_30 = b[30] ? a : 0;
assign pwire_31 = b[31] ? (~a) : 0;

endmodule